<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="swimrankings.net" version="5.77112">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Katowice" name="Puchar Polski Masters w Pływaniu" course="SCM" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2023-05-13" type="YEAR" />
      <POOL lanemin="1" lanemax="8" />
      <FACILITY city="Katowice" nation="POL" />
      <POINTTABLE pointtableid="3015" name="FINA Point Scoring" version="2022" />
      <SESSIONS>
        <SESSION date="2023-05-13" daytime="16:00" number="1">
          <EVENTS>
            <EVENT eventid="1" daytime="16:13" gender="M" number="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809836" />
                    <RANKING order="2" place="2" resultid="175810062" />
                    <RANKING order="3" place="3" resultid="175809896" />
                    <RANKING order="4" place="4" resultid="175810139" />
                    <RANKING order="5" place="5" resultid="175810351" />
                    <RANKING order="6" place="6" resultid="175810086" />
                    <RANKING order="7" place="7" resultid="175810518" />
                    <RANKING order="8" place="8" resultid="175810399" />
                    <RANKING order="9" place="9" resultid="175810024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810573" />
                    <RANKING order="2" place="2" resultid="175810133" />
                    <RANKING order="3" place="3" resultid="175810526" />
                    <RANKING order="4" place="4" resultid="175810458" />
                    <RANKING order="5" place="5" resultid="175809846" />
                    <RANKING order="6" place="6" resultid="175809991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810251" />
                    <RANKING order="2" place="2" resultid="175810300" />
                    <RANKING order="3" place="3" resultid="175810533" />
                    <RANKING order="4" place="4" resultid="175810563" />
                    <RANKING order="5" place="5" resultid="175810539" />
                    <RANKING order="6" place="6" resultid="175810093" />
                    <RANKING order="7" place="7" resultid="175810072" />
                    <RANKING order="8" place="8" resultid="175809852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810454" />
                    <RANKING order="2" place="2" resultid="175810577" />
                    <RANKING order="3" place="3" resultid="175809900" />
                    <RANKING order="4" place="4" resultid="175810137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810481" />
                    <RANKING order="2" place="2" resultid="175810017" />
                    <RANKING order="3" place="3" resultid="175810477" />
                    <RANKING order="4" place="4" resultid="175809920" />
                    <RANKING order="5" place="5" resultid="175809904" />
                    <RANKING order="6" place="6" resultid="175810547" />
                    <RANKING order="7" place="7" resultid="175809954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810261" />
                    <RANKING order="2" place="2" resultid="175810240" />
                    <RANKING order="3" place="3" resultid="175809932" />
                    <RANKING order="4" place="4" resultid="175810294" />
                    <RANKING order="5" place="5" resultid="175810290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810181" />
                    <RANKING order="2" place="2" resultid="175810084" />
                    <RANKING order="3" place="3" resultid="175809974" />
                    <RANKING order="4" place="4" resultid="175810354" />
                    <RANKING order="5" place="5" resultid="175810569" />
                    <RANKING order="6" place="6" resultid="175810189" />
                    <RANKING order="7" place="7" resultid="175810306" />
                    <RANKING order="8" place="8" resultid="175810417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809978" />
                    <RANKING order="2" place="2" resultid="175810395" />
                    <RANKING order="3" place="3" resultid="175810020" />
                    <RANKING order="4" place="4" resultid="175810099" />
                    <RANKING order="5" place="5" resultid="175810322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809994" />
                    <RANKING order="2" place="2" resultid="175810445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810460" />
                    <RANKING order="2" place="2" resultid="175810555" />
                    <RANKING order="3" place="3" resultid="175810043" />
                    <RANKING order="4" place="4" resultid="175810543" />
                    <RANKING order="5" place="5" resultid="175810268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810361" />
                    <RANKING order="2" place="2" resultid="175810607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="-1" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810377" />
                    <RANKING order="2" place="2" resultid="175810599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810333" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2" number="8" />
                <HEAT heatid="3" number="2" />
                <HEAT heatid="6" number="7" />
                <HEAT heatid="7" number="6" />
                <HEAT heatid="8" number="12" />
                <HEAT heatid="11" number="5" />
                <HEAT heatid="12" number="11" />
                <HEAT heatid="13" number="1" />
                <HEAT heatid="14" number="3" />
                <HEAT heatid="17" number="9" />
                <HEAT heatid="18" number="10" />
                <HEAT heatid="19" number="4" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2" daytime="16:00" gender="F" number="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810007" />
                    <RANKING order="2" place="2" resultid="175809873" />
                    <RANKING order="3" place="3" resultid="175810223" />
                    <RANKING order="4" place="4" resultid="175809966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810201" />
                    <RANKING order="2" place="2" resultid="175809983" />
                    <RANKING order="3" place="3" resultid="175810249" />
                    <RANKING order="4" place="4" resultid="175809940" />
                    <RANKING order="5" place="5" resultid="175809928" />
                    <RANKING order="6" place="6" resultid="175810068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810465" />
                    <RANKING order="2" place="2" resultid="175810177" />
                    <RANKING order="3" place="3" resultid="175810565" />
                    <RANKING order="4" place="4" resultid="175809958" />
                    <RANKING order="5" place="5" resultid="175810385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810047" />
                    <RANKING order="2" place="2" resultid="175810153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="-1" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810060" />
                    <RANKING order="2" place="2" resultid="175810070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810149" />
                    <RANKING order="2" place="2" resultid="175810286" />
                    <RANKING order="3" place="3" resultid="175810296" />
                    <RANKING order="4" place="4" resultid="175810065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810318" />
                    <RANKING order="2" place="2" resultid="175810081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810522" />
                    <RANKING order="2" place="2" resultid="175810331" />
                    <RANKING order="3" place="3" resultid="175810347" />
                    <RANKING order="4" place="4" resultid="175810244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810389" />
                    <RANKING order="2" place="2" resultid="175810365" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4" number="5" />
                <HEAT heatid="5" number="4" />
                <HEAT heatid="9" number="3" />
                <HEAT heatid="10" number="1" />
                <HEAT heatid="15" number="6" />
                <HEAT heatid="16" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5" daytime="17:49" gender="M" number="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809837" />
                    <RANKING order="2" place="2" resultid="175810370" />
                    <RANKING order="3" place="3" resultid="175810140" />
                    <RANKING order="4" place="4" resultid="175810519" />
                    <RANKING order="5" place="5" resultid="175810025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810134" />
                    <RANKING order="2" place="2" resultid="175810574" />
                    <RANKING order="3" place="3" resultid="175810170" />
                    <RANKING order="4" place="4" resultid="175810107" />
                    <RANKING order="5" place="5" resultid="175810459" />
                    <RANKING order="6" place="6" resultid="175809847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809962" />
                    <RANKING order="2" place="2" resultid="175810216" />
                    <RANKING order="3" place="3" resultid="175810021" />
                    <RANKING order="4" place="4" resultid="175810396" />
                    <RANKING order="5" place="5" resultid="175810100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810161" />
                    <RANKING order="2" place="2" resultid="175810257" />
                    <RANKING order="3" place="3" resultid="175810570" />
                    <RANKING order="4" place="4" resultid="175810355" />
                    <RANKING order="5" place="5" resultid="175810307" />
                    <RANKING order="6" place="6" resultid="175810245" />
                    <RANKING order="7" place="7" resultid="175810190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810578" />
                    <RANKING order="2" place="2" resultid="175810174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810581" />
                    <RANKING order="2" place="2" resultid="175810381" />
                    <RANKING order="3" place="3" resultid="175810337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810378" />
                    <RANKING order="2" place="2" resultid="175810600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810604" />
                    <RANKING order="2" place="2" resultid="175810608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810544" />
                    <RANKING order="2" place="2" resultid="175810233" />
                    <RANKING order="3" place="3" resultid="175810269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810334" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="35" number="5" />
                <HEAT heatid="36" number="1" />
                <HEAT heatid="39" number="7" />
                <HEAT heatid="40" number="2" />
                <HEAT heatid="42" number="6" />
                <HEAT heatid="43" number="4" />
                <HEAT heatid="44" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6" daytime="17:27" gender="F" number="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810178" />
                    <RANKING order="2" place="2" resultid="175809860" />
                    <RANKING order="3" place="3" resultid="175810466" />
                    <RANKING order="4" place="4" resultid="175810566" />
                    <RANKING order="5" place="5" resultid="175810473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810451" />
                    <RANKING order="2" place="2" resultid="175810042" />
                    <RANKING order="3" place="3" resultid="175809941" />
                    <RANKING order="4" place="4" resultid="175810314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810048" />
                    <RANKING order="2" place="2" resultid="175810255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810492" />
                    <RANKING order="2" place="2" resultid="175810287" />
                    <RANKING order="3" place="3" resultid="175810066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810374" />
                    <RANKING order="2" place="2" resultid="175810231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810502" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="37" number="4" />
                <HEAT heatid="38" number="2" />
                <HEAT heatid="41" number="1" />
                <HEAT heatid="45" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="11" daytime="16:45" gender="M" number="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809970" />
                    <RANKING order="2" place="2" resultid="175810212" />
                    <RANKING order="3" place="3" resultid="175810235" />
                    <RANKING order="4" place="4" resultid="175810089" />
                    <RANKING order="5" place="5" resultid="175809856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810343" />
                    <RANKING order="2" place="2" resultid="175809866" />
                    <RANKING order="3" place="3" resultid="175810369" />
                    <RANKING order="4" place="4" resultid="175810400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809881" />
                    <RANKING order="2" place="2" resultid="175810279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810165" />
                    <RANKING order="2" place="2" resultid="175810169" />
                    <RANKING order="3" place="3" resultid="175810111" />
                    <RANKING order="4" place="4" resultid="175809892" />
                    <RANKING order="5" place="5" resultid="175810562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809921" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810129" />
                    <RANKING order="2" place="2" resultid="175810078" />
                    <RANKING order="3" place="3" resultid="175810103" />
                    <RANKING order="4" place="4" resultid="175810256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810119" />
                    <RANKING order="2" place="2" resultid="175810506" />
                    <RANKING order="3" place="3" resultid="175810603" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810228" />
                    <RANKING order="2" place="2" resultid="175810173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810193" />
                    <RANKING order="2" place="2" resultid="175810252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810499" />
                    <RANKING order="2" place="2" resultid="175810446" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="63" number="2" />
                <HEAT heatid="64" number="3" />
                <HEAT heatid="66" number="1" />
                <HEAT heatid="67" number="4" />
                <HEAT heatid="70" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="12" daytime="16:34" gender="F" number="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809874" />
                    <RANKING order="2" place="2" resultid="175810437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809984" />
                    <RANKING order="2" place="2" resultid="175810041" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810220" />
                    <RANKING order="2" place="2" resultid="175810001" />
                    <RANKING order="3" place="3" resultid="175810283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810441" />
                    <RANKING order="2" place="2" resultid="175810028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810405" />
                    <RANKING order="2" place="2" resultid="175810595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810491" />
                    <RANKING order="2" place="2" resultid="175810297" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="65" number="3" />
                <HEAT heatid="68" number="1" />
                <HEAT heatid="69" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="15" daytime="16:59" gender="F" number="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810202" />
                    <RANKING order="2" place="2" resultid="175809929" />
                    <RANKING order="3" place="3" resultid="175809916" />
                    <RANKING order="4" place="4" resultid="175809840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809924" />
                    <RANKING order="2" place="2" resultid="175810208" />
                    <RANKING order="3" place="3" resultid="175809843" />
                    <RANKING order="4" place="-1" resultid="175809913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809863" />
                    <RANKING order="2" place="2" resultid="175810057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810185" />
                    <RANKING order="2" place="2" resultid="175810074" />
                    <RANKING order="3" place="3" resultid="175809959" />
                    <RANKING order="4" place="4" resultid="175810386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810008" />
                    <RANKING order="2" place="2" resultid="175810224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810591" />
                    <RANKING order="2" place="2" resultid="175810121" />
                    <RANKING order="3" place="3" resultid="175810051" />
                    <RANKING order="4" place="4" resultid="175810011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810145" />
                    <RANKING order="2" place="2" resultid="175810449" />
                    <RANKING order="3" place="3" resultid="175810082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810523" />
                    <RANKING order="2" place="2" resultid="175810327" />
                    <RANKING order="3" place="3" resultid="175810514" />
                    <RANKING order="4" place="4" resultid="175810243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810430" />
                    <RANKING order="2" place="2" resultid="175810366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810413" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="77" number="1" />
                <HEAT heatid="78" number="2" />
                <HEAT heatid="80" number="5" />
                <HEAT heatid="85" number="4" />
                <HEAT heatid="86" number="3" />
                <HEAT heatid="88" number="6" />
              </HEATS>
            </EVENT>
            <EVENT eventid="16" daytime="17:11" gender="M" number="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810585" />
                    <RANKING order="2" place="2" resultid="175809884" />
                    <RANKING order="3" place="3" resultid="175809857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809867" />
                    <RANKING order="2" place="2" resultid="175810037" />
                    <RANKING order="3" place="3" resultid="175810087" />
                    <RANKING order="4" place="4" resultid="175810265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810125" />
                    <RANKING order="2" place="2" resultid="175810073" />
                    <RANKING order="3" place="3" resultid="175809877" />
                    <RANKING order="4" place="4" resultid="175810540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809888" />
                    <RANKING order="2" place="2" resultid="175810464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810018" />
                    <RANKING order="2" place="2" resultid="175810271" />
                    <RANKING order="3" place="3" resultid="175809905" />
                    <RANKING order="4" place="4" resultid="175810469" />
                    <RANKING order="5" place="5" resultid="175810548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810182" />
                    <RANKING order="2" place="2" resultid="175809982" />
                    <RANKING order="3" place="3" resultid="175810403" />
                    <RANKING order="4" place="4" resultid="175809975" />
                    <RANKING order="5" place="5" resultid="175809908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810262" />
                    <RANKING order="2" place="2" resultid="175810495" />
                    <RANKING order="3" place="3" resultid="175810275" />
                    <RANKING order="4" place="4" resultid="175810295" />
                    <RANKING order="5" place="5" resultid="175809933" />
                    <RANKING order="6" place="6" resultid="175810529" />
                    <RANKING order="7" place="7" resultid="175810291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810055" />
                    <RANKING order="2" place="2" resultid="175810427" />
                    <RANKING order="3" place="3" resultid="175810138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810115" />
                    <RANKING order="2" place="2" resultid="175810310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810424" />
                    <RANKING order="2" place="2" resultid="175810157" />
                    <RANKING order="3" place="3" resultid="175810535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810362" />
                    <RANKING order="2" place="2" resultid="175810559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="-1" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810510" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="79" number="3" />
                <HEAT heatid="81" number="1" />
                <HEAT heatid="82" number="4" />
                <HEAT heatid="83" number="5" />
                <HEAT heatid="84" number="7" />
                <HEAT heatid="87" number="6" />
                <HEAT heatid="89" number="8" />
                <HEAT heatid="90" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19" daytime="19:06" gender="F" number="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809917" />
                    <RANKING order="2" place="2" resultid="175809841" />
                    <RANKING order="3" place="3" resultid="175810069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810392" />
                    <RANKING order="2" place="2" resultid="175809925" />
                    <RANKING order="3" place="3" resultid="175809945" />
                    <RANKING order="4" place="4" resultid="175809844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810592" />
                    <RANKING order="2" place="2" resultid="175810012" />
                    <RANKING order="3" place="3" resultid="175810052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810058" />
                    <RANKING order="2" place="2" resultid="175810410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810186" />
                    <RANKING order="2" place="2" resultid="175810075" />
                    <RANKING order="3" place="3" resultid="175810421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810146" />
                    <RANKING order="2" place="2" resultid="175810450" />
                    <RANKING order="3" place="3" resultid="175810083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810431" />
                    <RANKING order="2" place="2" resultid="175810232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810414" />
                    <RANKING order="2" place="2" resultid="175810340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810503" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="102" number="1" />
                <HEAT heatid="108" number="3" />
                <HEAT heatid="109" number="4" />
                <HEAT heatid="111" number="2" />
                <HEAT heatid="112" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="20" daytime="19:40" gender="M" number="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810126" />
                    <RANKING order="2" place="2" resultid="175810301" />
                    <RANKING order="3" place="3" resultid="175809878" />
                    <RANKING order="4" place="4" resultid="175809853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810158" />
                    <RANKING order="2" place="2" resultid="175810425" />
                    <RANKING order="3" place="3" resultid="175809882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810586" />
                    <RANKING order="2" place="2" resultid="175809971" />
                    <RANKING order="3" place="3" resultid="175809885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810162" />
                    <RANKING order="2" place="2" resultid="175810104" />
                    <RANKING order="3" place="3" resultid="175809909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810056" />
                    <RANKING order="2" place="2" resultid="175810428" />
                    <RANKING order="3" place="3" resultid="175810014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810112" />
                    <RANKING order="2" place="2" resultid="175810116" />
                    <RANKING order="3" place="3" resultid="175810108" />
                    <RANKING order="4" place="4" resultid="175810311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810344" />
                    <RANKING order="2" place="2" resultid="175810266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810496" />
                    <RANKING order="2" place="2" resultid="175810276" />
                    <RANKING order="3" place="3" resultid="175810530" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="103" number="1" />
                <HEAT heatid="104" number="2" />
                <HEAT heatid="105" number="6" />
                <HEAT heatid="106" number="3" />
                <HEAT heatid="107" number="4" />
                <HEAT heatid="110" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="23" daytime="18:52" gender="F" number="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809861" />
                    <RANKING order="2" place="2" resultid="175810474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810319" />
                    <RANKING order="2" place="2" resultid="175809937" />
                    <RANKING order="3" place="3" resultid="175810002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809988" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="123" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="24" daytime="18:55" gender="M" number="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810482" />
                    <RANKING order="2" place="2" resultid="175810272" />
                    <RANKING order="3" place="3" resultid="175810478" />
                    <RANKING order="4" place="4" resultid="175809955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809963" />
                    <RANKING order="2" place="2" resultid="175810213" />
                    <RANKING order="3" place="3" resultid="175809979" />
                    <RANKING order="4" place="4" resultid="175810090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810455" />
                    <RANKING order="2" place="2" resultid="175810013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810085" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810582" />
                    <RANKING order="2" place="2" resultid="175810382" />
                    <RANKING order="3" place="3" resultid="175810239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810461" />
                    <RANKING order="2" place="2" resultid="175810280" />
                    <RANKING order="3" place="3" resultid="175810234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810507" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="124" number="2" />
                <HEAT heatid="125" number="4" />
                <HEAT heatid="126" number="3" />
                <HEAT heatid="127" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="27" daytime="18:20" gender="F" number="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809870" />
                    <RANKING order="2" place="2" resultid="175809936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809944" />
                    <RANKING order="2" place="2" resultid="175809998" />
                    <RANKING order="3" place="-1" resultid="175810391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810444" />
                    <RANKING order="2" place="2" resultid="175810409" />
                    <RANKING order="3" place="3" resultid="175810029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810150" />
                    <RANKING order="2" place="2" resultid="175810122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810406" />
                    <RANKING order="2" place="2" resultid="175810596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810328" />
                    <RANKING order="2" place="2" resultid="175810515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810316" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="131" number="3" />
                <HEAT heatid="134" number="1" />
                <HEAT heatid="135" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="28" daytime="18:37" gender="M" number="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809897" />
                    <RANKING order="2" place="2" resultid="175810088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810536" />
                    <RANKING order="2" place="2" resultid="175810556" />
                    <RANKING order="3" place="3" resultid="175810044" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810130" />
                    <RANKING order="2" place="2" resultid="175810246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810194" />
                    <RANKING order="2" place="2" resultid="175810564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810217" />
                    <RANKING order="2" place="2" resultid="175810236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810260" />
                    <RANKING order="2" place="2" resultid="175810470" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="132" number="2" />
                <HEAT heatid="133" number="1" />
                <HEAT heatid="136" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="31" daytime="20:09" gender="X" number="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="199" agemin="160">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810199" />
                    <RANKING order="2" place="2" resultid="175809952" />
                    <RANKING order="3" place="3" resultid="175810325" />
                    <RANKING order="4" place="4" resultid="175809850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="279" agemin="240">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809948" />
                    <RANKING order="2" place="2" resultid="175810032" />
                    <RANKING order="3" place="3" resultid="175810418" />
                    <RANKING order="4" place="4" resultid="175810034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="239" agemin="200">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810036" />
                    <RANKING order="2" place="2" resultid="175809950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="159" agemin="120">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810197" />
                    <RANKING order="2" place="2" resultid="175810304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="119" agemin="100">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810485" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="148" number="2" />
                <HEAT heatid="149" number="3" />
                <HEAT heatid="150" number="1" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2023-05-14" daytime="08:45" number="2">
          <EVENTS>
            <EVENT eventid="3" daytime="09:32" gender="M" number="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809838" />
                    <RANKING order="2" place="2" resultid="175810345" />
                    <RANKING order="3" place="3" resultid="175810141" />
                    <RANKING order="4" place="4" resultid="175810401" />
                    <RANKING order="5" place="5" resultid="175810026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810117" />
                    <RANKING order="2" place="2" resultid="175810575" />
                    <RANKING order="3" place="3" resultid="175810135" />
                    <RANKING order="4" place="4" resultid="175810171" />
                    <RANKING order="5" place="5" resultid="175810527" />
                    <RANKING order="6" place="6" resultid="175810109" />
                    <RANKING order="7" place="7" resultid="175809894" />
                    <RANKING order="8" place="8" resultid="175809848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810218" />
                    <RANKING order="2" place="2" resultid="175810397" />
                    <RANKING order="3" place="3" resultid="175809886" />
                    <RANKING order="4" place="4" resultid="175810237" />
                    <RANKING order="5" place="5" resultid="175810323" />
                    <RANKING order="6" place="6" resultid="175810206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810456" />
                    <RANKING order="2" place="2" resultid="175810580" />
                    <RANKING order="3" place="3" resultid="175809902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810583" />
                    <RANKING order="2" place="2" resultid="175810383" />
                    <RANKING order="3" place="3" resultid="175810497" />
                    <RANKING order="4" place="4" resultid="175809934" />
                    <RANKING order="5" place="5" resultid="175810487" />
                    <RANKING order="6" place="6" resultid="175810292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809976" />
                    <RANKING order="2" place="2" resultid="175810356" />
                    <RANKING order="3" place="3" resultid="175810005" />
                    <RANKING order="4" place="4" resultid="175810572" />
                    <RANKING order="5" place="5" resultid="175810191" />
                    <RANKING order="6" place="6" resultid="175810308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809996" />
                    <RANKING order="2" place="2" resultid="175810447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810097" />
                    <RANKING order="2" place="2" resultid="175810019" />
                    <RANKING order="3" place="3" resultid="175810484" />
                    <RANKING order="4" place="4" resultid="175810471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810552" />
                    <RANKING order="2" place="2" resultid="175810144" />
                    <RANKING order="3" place="3" resultid="175810534" />
                    <RANKING order="4" place="4" resultid="175810541" />
                    <RANKING order="5" place="5" resultid="175810095" />
                    <RANKING order="6" place="6" resultid="175810207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810462" />
                    <RANKING order="2" place="2" resultid="175810557" />
                    <RANKING order="3" place="3" resultid="175810537" />
                    <RANKING order="4" place="4" resultid="175810545" />
                    <RANKING order="5" place="5" resultid="175810270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810380" />
                    <RANKING order="2" place="2" resultid="175810601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810605" />
                    <RANKING order="2" place="2" resultid="175810609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810336" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20" number="8" />
                <HEAT heatid="21" number="2" />
                <HEAT heatid="24" number="6" />
                <HEAT heatid="25" number="5" />
                <HEAT heatid="28" number="7" />
                <HEAT heatid="29" number="4" />
                <HEAT heatid="30" number="11" />
                <HEAT heatid="31" number="3" />
                <HEAT heatid="32" number="1" />
                <HEAT heatid="33" number="10" />
                <HEAT heatid="34" number="9" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4" daytime="09:17" gender="F" number="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809864" />
                    <RANKING order="2" place="2" resultid="175809989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809875" />
                    <RANKING order="2" place="2" resultid="175810225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810452" />
                    <RANKING order="2" place="2" resultid="175810204" />
                    <RANKING order="3" place="3" resultid="175810250" />
                    <RANKING order="4" place="4" resultid="175809943" />
                    <RANKING order="5" place="5" resultid="175809930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810179" />
                    <RANKING order="2" place="2" resultid="175810467" />
                    <RANKING order="3" place="3" resultid="175810568" />
                    <RANKING order="4" place="4" resultid="175809960" />
                    <RANKING order="5" place="5" resultid="175810387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810288" />
                    <RANKING order="2" place="2" resultid="175810067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810504" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="22" number="3" />
                <HEAT heatid="23" number="4" />
                <HEAT heatid="26" number="2" />
                <HEAT heatid="27" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7" daytime="12:46" gender="M" number="32" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810136" />
                    <RANKING order="2" place="2" resultid="175810118" />
                    <RANKING order="3" place="3" resultid="175810490" />
                    <RANKING order="4" place="4" resultid="175810110" />
                    <RANKING order="5" place="5" resultid="175809895" />
                    <RANKING order="6" place="6" resultid="175809849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809965" />
                    <RANKING order="2" place="2" resultid="175810219" />
                    <RANKING order="3" place="3" resultid="175810238" />
                    <RANKING order="4" place="4" resultid="175809887" />
                    <RANKING order="5" place="5" resultid="175810092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810132" />
                    <RANKING order="2" place="2" resultid="175810164" />
                    <RANKING order="3" place="3" resultid="175810006" />
                    <RANKING order="4" place="4" resultid="175810259" />
                    <RANKING order="5" place="5" resultid="175810248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810372" />
                    <RANKING order="2" place="2" resultid="175810521" />
                    <RANKING order="3" place="3" resultid="175810027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810160" />
                    <RANKING order="2" place="2" resultid="175810546" />
                    <RANKING order="3" place="3" resultid="175810282" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810584" />
                    <RANKING order="2" place="2" resultid="175810488" />
                    <RANKING order="3" place="3" resultid="175810338" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="46" number="2" />
                <HEAT heatid="47" number="4" />
                <HEAT heatid="48" number="5" />
                <HEAT heatid="50" number="1" />
                <HEAT heatid="52" number="6" />
                <HEAT heatid="54" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8" daytime="12:14" gender="F" number="31" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810443" />
                    <RANKING order="2" place="2" resultid="175810031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810453" />
                    <RANKING order="2" place="2" resultid="175810315" />
                    <RANKING order="3" place="3" resultid="175810554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810598" />
                    <RANKING order="2" place="2" resultid="175810342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810505" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="49" number="2" />
                <HEAT heatid="51" number="1" />
                <HEAT heatid="53" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="9" daytime="12:04" gender="M" number="30" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809839" />
                    <RANKING order="2" place="2" resultid="175809869" />
                    <RANKING order="3" place="3" resultid="175810142" />
                    <RANKING order="4" place="4" resultid="175810353" />
                    <RANKING order="5" place="5" resultid="175810402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810023" />
                    <RANKING order="2" place="2" resultid="175810324" />
                    <RANKING order="3" place="3" resultid="175809859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810098" />
                    <RANKING order="2" place="2" resultid="175809907" />
                    <RANKING order="3" place="3" resultid="175810480" />
                    <RANKING order="4" place="4" resultid="175810550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810168" />
                    <RANKING order="2" place="2" resultid="175810528" />
                    <RANKING order="3" place="3" resultid="175809993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810080" />
                    <RANKING order="2" place="2" resultid="175810106" />
                    <RANKING order="3" place="3" resultid="175810309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810254" />
                    <RANKING order="2" place="2" resultid="175810196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810501" />
                    <RANKING order="2" place="2" resultid="175810448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810513" />
                    <RANKING order="2" place="2" resultid="175810602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810509" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="55" number="4" />
                <HEAT heatid="56" number="2" />
                <HEAT heatid="57" number="3" />
                <HEAT heatid="59" number="5" />
                <HEAT heatid="60" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10" daytime="11:55" gender="F" number="29" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809876" />
                    <RANKING order="2" place="2" resultid="175810227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809986" />
                    <RANKING order="2" place="2" resultid="175810590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810222" />
                    <RANKING order="2" place="2" resultid="175810004" />
                    <RANKING order="3" place="3" resultid="175810285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810152" />
                    <RANKING order="2" place="2" resultid="175810494" />
                    <RANKING order="3" place="3" resultid="175810299" />
                    <RANKING order="4" place="4" resultid="175810054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810061" />
                    <RANKING order="2" place="2" resultid="175810071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810423" />
                    <RANKING order="2" place="2" resultid="175810388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810416" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="58" number="3" />
                <HEAT heatid="61" number="2" />
                <HEAT heatid="62" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="13" daytime="10:52" gender="M" number="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809973" />
                    <RANKING order="2" place="2" resultid="175810091" />
                    <RANKING order="3" place="3" resultid="175809858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810079" />
                    <RANKING order="2" place="2" resultid="175810258" />
                    <RANKING order="3" place="3" resultid="175810247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810120" />
                    <RANKING order="2" place="2" resultid="175810508" />
                    <RANKING order="3" place="3" resultid="175810606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810229" />
                    <RANKING order="2" place="2" resultid="175810175" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810195" />
                    <RANKING order="2" place="2" resultid="175810253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810371" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="71" number="2" />
                <HEAT heatid="73" number="3" />
                <HEAT heatid="75" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="14" daytime="10:34" gender="F" number="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810221" />
                    <RANKING order="2" place="2" resultid="175810284" />
                    <RANKING order="3" place="3" resultid="175809938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809985" />
                    <RANKING order="2" place="2" resultid="175810553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810597" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="72" number="3" />
                <HEAT heatid="74" number="2" />
                <HEAT heatid="76" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="17" daytime="10:00" gender="F" number="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810589" />
                    <RANKING order="2" place="2" resultid="175809919" />
                    <RANKING order="3" place="3" resultid="175809842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810393" />
                    <RANKING order="2" place="2" resultid="175809926" />
                    <RANKING order="3" place="3" resultid="175810209" />
                    <RANKING order="4" place="4" resultid="175809915" />
                    <RANKING order="5" place="5" resultid="175809845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810187" />
                    <RANKING order="2" place="2" resultid="175810076" />
                    <RANKING order="3" place="3" resultid="175809961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810593" />
                    <RANKING order="2" place="2" resultid="175810053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810059" />
                    <RANKING order="2" place="2" resultid="175810411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810359" />
                    <RANKING order="2" place="2" resultid="175810147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810433" />
                    <RANKING order="2" place="2" resultid="175810367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810415" />
                    <RANKING order="2" place="2" resultid="175810341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810329" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="91" number="2" />
                <HEAT heatid="92" number="1" />
                <HEAT heatid="97" number="3" />
                <HEAT heatid="98" number="4" />
                <HEAT heatid="101" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="18" daytime="10:17" gender="M" number="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810542" />
                    <RANKING order="2" place="2" resultid="175809879" />
                    <RANKING order="3" place="3" resultid="175809854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809868" />
                    <RANKING order="2" place="2" resultid="175810039" />
                    <RANKING order="3" place="3" resultid="175810267" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810426" />
                    <RANKING order="2" place="2" resultid="175810159" />
                    <RANKING order="3" place="3" resultid="175809883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810274" />
                    <RANKING order="2" place="2" resultid="175809906" />
                    <RANKING order="3" place="3" resultid="175810549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810587" />
                    <RANKING order="2" place="2" resultid="175809972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810429" />
                    <RANKING order="2" place="2" resultid="175810015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810183" />
                    <RANKING order="2" place="2" resultid="175810105" />
                    <RANKING order="3" place="3" resultid="175810404" />
                    <RANKING order="4" place="-1" resultid="175810357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810113" />
                    <RANKING order="2" place="2" resultid="175810312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810263" />
                    <RANKING order="2" place="2" resultid="175810498" />
                    <RANKING order="3" place="3" resultid="175810278" />
                    <RANKING order="4" place="4" resultid="175810531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="-1" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810561" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="93" number="1" />
                <HEAT heatid="94" number="3" />
                <HEAT heatid="95" number="6" />
                <HEAT heatid="96" number="5" />
                <HEAT heatid="99" number="4" />
                <HEAT heatid="100" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="21" daytime="08:57" gender="F" number="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809871" />
                    <RANKING order="2" place="2" resultid="175810003" />
                    <RANKING order="3" place="3" resultid="175810320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810203" />
                    <RANKING order="2" place="2" resultid="175809942" />
                    <RANKING order="3" place="3" resultid="175809918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810009" />
                    <RANKING order="2" place="2" resultid="175809968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810524" />
                    <RANKING order="2" place="2" resultid="175810516" />
                    <RANKING order="3" place="3" resultid="175810349" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="113" number="3" />
                <HEAT heatid="116" number="1" />
                <HEAT heatid="118" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="22" daytime="09:04" gender="M" number="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809898" />
                    <RANKING order="2" place="2" resultid="175810063" />
                    <RANKING order="3" place="3" resultid="175810352" />
                    <RANKING order="4" place="4" resultid="175810038" />
                    <RANKING order="5" place="5" resultid="175810520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809910" />
                    <RANKING order="2" place="2" resultid="175810571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810483" />
                    <RANKING order="2" place="2" resultid="175810479" />
                    <RANKING order="3" place="3" resultid="175809922" />
                    <RANKING order="4" place="4" resultid="175810273" />
                    <RANKING order="5" place="5" resultid="175809956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809980" />
                    <RANKING order="2" place="2" resultid="175810214" />
                    <RANKING order="3" place="3" resultid="175810022" />
                    <RANKING order="4" place="4" resultid="175810101" />
                    <RANKING order="5" place="5" resultid="175810205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810045" />
                    <RANKING order="2" place="2" resultid="175810281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810551" />
                    <RANKING order="2" place="2" resultid="175810127" />
                    <RANKING order="3" place="3" resultid="175810143" />
                    <RANKING order="4" place="4" resultid="175810302" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810241" />
                    <RANKING order="2" place="2" resultid="175810532" />
                    <RANKING order="3" place="3" resultid="175810277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="-1" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810379" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="114" number="5" />
                <HEAT heatid="115" number="3" />
                <HEAT heatid="117" number="7" />
                <HEAT heatid="119" number="4" />
                <HEAT heatid="120" number="6" />
                <HEAT heatid="121" number="2" />
                <HEAT heatid="122" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="25" daytime="11:13" gender="M" number="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810163" />
                    <RANKING order="2" place="2" resultid="175809911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809964" />
                    <RANKING order="2" place="2" resultid="175810215" />
                    <RANKING order="3" place="3" resultid="175810102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810489" />
                    <RANKING order="2" place="2" resultid="175810114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810463" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="128" number="2" />
                <HEAT heatid="130" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="26" daytime="11:07" gender="F" number="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809990" />
                    <RANKING order="2" place="2" resultid="175810412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810124" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810475" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="129" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="29" daytime="11:24" gender="F" number="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809865" />
                    <RANKING order="2" place="2" resultid="175810030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809872" />
                    <RANKING order="2" place="2" resultid="175810148" />
                    <RANKING order="3" place="3" resultid="175810321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810394" />
                    <RANKING order="2" place="2" resultid="175809927" />
                    <RANKING order="3" place="3" resultid="175810210" />
                    <RANKING order="4" place="4" resultid="175810000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810317" />
                    <RANKING order="2" place="2" resultid="175809931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810010" />
                    <RANKING order="2" place="2" resultid="175809969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810180" />
                    <RANKING order="2" place="2" resultid="175810468" />
                    <RANKING order="3" place="3" resultid="175810188" />
                    <RANKING order="4" place="4" resultid="175810077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810151" />
                    <RANKING order="2" place="2" resultid="175810594" />
                    <RANKING order="3" place="3" resultid="175810298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810330" />
                    <RANKING order="2" place="2" resultid="175810525" />
                    <RANKING order="3" place="3" resultid="175810517" />
                    <RANKING order="4" place="4" resultid="175810350" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="137" number="3" />
                <HEAT heatid="138" number="4" />
                <HEAT heatid="143" number="2" />
                <HEAT heatid="145" number="1" />
                <HEAT heatid="146" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="30" daytime="11:39" gender="M" number="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810303" />
                    <RANKING order="2" place="2" resultid="175809880" />
                    <RANKING order="3" place="3" resultid="175810096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810346" />
                    <RANKING order="2" place="2" resultid="175809899" />
                    <RANKING order="3" place="3" resultid="175810064" />
                    <RANKING order="4" place="4" resultid="175810040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810457" />
                    <RANKING order="2" place="-1" resultid="175809903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809923" />
                    <RANKING order="2" place="2" resultid="175810472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810264" />
                    <RANKING order="2" place="2" resultid="175810242" />
                    <RANKING order="3" place="3" resultid="175809935" />
                    <RANKING order="4" place="4" resultid="175810293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810131" />
                    <RANKING order="2" place="2" resultid="175810184" />
                    <RANKING order="3" place="3" resultid="175809977" />
                    <RANKING order="4" place="4" resultid="175810192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810588" />
                    <RANKING order="2" place="2" resultid="175809981" />
                    <RANKING order="3" place="3" resultid="175810398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810172" />
                    <RANKING order="2" place="2" resultid="175810576" />
                    <RANKING order="3" place="3" resultid="175810313" />
                    <RANKING order="4" place="4" resultid="175809992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810558" />
                    <RANKING order="2" place="2" resultid="175810538" />
                    <RANKING order="3" place="3" resultid="175810046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810364" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="139" number="2" />
                <HEAT heatid="140" number="1" />
                <HEAT heatid="141" number="3" />
                <HEAT heatid="142" number="6" />
                <HEAT heatid="144" number="4" />
                <HEAT heatid="147" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="32" daytime="08:45" gender="X" number="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="199" agemin="160">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809953" />
                    <RANKING order="2" place="2" resultid="175810326" />
                    <RANKING order="3" place="3" resultid="175810211" />
                    <RANKING order="4" place="4" resultid="175809851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="279" agemin="240">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175809949" />
                    <RANKING order="2" place="2" resultid="175810033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="239" agemin="200">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810200" />
                    <RANKING order="2" place="2" resultid="175810035" />
                    <RANKING order="3" place="3" resultid="175809951" />
                    <RANKING order="4" place="4" resultid="175810419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="159" agemin="120">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810198" />
                    <RANKING order="2" place="2" resultid="175810305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="119" agemin="100">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="175810486" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="151" number="2" />
                <HEAT heatid="152" number="1" />
                <HEAT heatid="153" number="3" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="POL" region="UNT" clubid="75947" swrid="75947" name="Start Katowice">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Slosarczyk" birthdate="1998-09-13" gender="M" nation="POL" swrid="5567825" athleteid="5567825">
              <HANDICAP breast="21" free="21" medley="21" />
              <RESULTS>
                <RESULT eventid="1" points="179" swimtime="00:00:35.77" resultid="175809954" heatid="11" lane="5" />
                <RESULT eventid="7" points="144" swimtime="00:06:44.05" resultid="175809957" heatid="47" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.35" />
                    <SPLIT distance="100" swimtime="00:01:34.09" />
                    <SPLIT distance="150" swimtime="00:02:27.11" />
                    <SPLIT distance="200" swimtime="00:03:20.57" />
                    <SPLIT distance="250" swimtime="00:04:13.70" />
                    <SPLIT distance="300" swimtime="00:05:05.80" />
                    <SPLIT distance="350" swimtime="00:05:57.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="160" swimtime="00:00:40.05" resultid="175809956" heatid="119" lane="5" />
                <RESULT eventid="24" points="125" swimtime="00:01:35.52" resultid="175809955" heatid="124" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03311" nation="POL" region="11" clubid="84349" swrid="84349" name="UKS Wodnik-29 Katowice" shortname="UKS Wodnik Katowice">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Korus" birthdate="1992-01-13" gender="M" nation="POL" swrid="4099337" athleteid="4099337">
              <RESULTS>
                <RESULT eventid="1" points="364" swimtime="00:00:28.23" resultid="175810043" heatid="2" lane="3" />
                <RESULT eventid="22" points="339" swimtime="00:00:31.19" resultid="175810045" heatid="114" lane="3" />
                <RESULT eventid="28" points="281" swimtime="00:02:47.27" resultid="175810044" heatid="132" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:16.76" />
                    <SPLIT distance="150" swimtime="00:02:06.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="302" swimtime="00:01:13.39" resultid="175810046" heatid="144" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Gawełczyk" birthdate="1991-07-26" gender="F" nation="POL" swrid="4072320" athleteid="4072320">
              <RESULTS>
                <RESULT eventid="2" points="542" swimtime="00:00:28.11" resultid="175810047" heatid="15" lane="5" />
                <RESULT eventid="6" points="533" swimtime="00:02:15.97" resultid="175810048" heatid="37" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:05.04" />
                    <SPLIT distance="150" swimtime="00:01:40.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" points="472" swimtime="00:00:31.30" resultid="175810049" heatid="113" lane="3" />
                <RESULT eventid="29" points="471" swimtime="00:01:12.61" resultid="175810050" heatid="146" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystyna" lastname="Nicpon" birthdate="1940-07-09" gender="F" nation="POL" swrid="4877349" athleteid="4877349">
              <RESULTS>
                <RESULT eventid="2" points="24" swimtime="00:01:18.83" resultid="175810060" heatid="16" lane="6" />
                <RESULT eventid="10" points="30" swimtime="00:01:21.21" resultid="175810061" heatid="61" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Wilczek" birthdate="1958-03-01" gender="M" nation="POL" swrid="4992641" athleteid="4992641">
              <RESULTS>
                <RESULT eventid="1" points="255" swimtime="00:00:31.79" resultid="175810062" heatid="2" lane="4" />
                <RESULT eventid="22" points="237" swimtime="00:00:35.13" resultid="175810063" heatid="114" lane="6" />
                <RESULT eventid="30" points="160" swimtime="00:01:30.63" resultid="175810064" heatid="141" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Głowacka" birthdate="1987-06-20" gender="F" nation="POL" swrid="5626905" athleteid="5626905">
              <RESULTS>
                <RESULT eventid="2" points="166" swimtime="00:00:41.65" resultid="175810065" heatid="9" lane="5" />
                <RESULT eventid="4" points="134" swimtime="00:01:37.97" resultid="175810067" heatid="26" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" points="123" swimtime="00:03:41.43" resultid="175810066" heatid="38" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.47" />
                    <SPLIT distance="100" swimtime="00:01:46.80" />
                    <SPLIT distance="150" swimtime="00:02:45.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Cichecka" birthdate="1982-01-01" gender="F" nation="POL" swrid="5626898" athleteid="5626898">
              <RESULTS>
                <RESULT eventid="2" points="171" swimtime="00:00:41.28" resultid="175810068" heatid="9" lane="6" />
                <RESULT eventid="19" points="97" swimtime="00:04:52.01" resultid="175810069" heatid="111" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.99" />
                    <SPLIT distance="100" swimtime="00:02:21.25" />
                    <SPLIT distance="150" swimtime="00:03:36.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Sieroń" birthdate="1981-01-01" gender="M" nation="POL" swrid="5626934" athleteid="5626934">
              <RESULTS>
                <RESULT eventid="1" points="177" swimtime="00:00:35.85" resultid="175810072" heatid="17" lane="2" />
                <RESULT eventid="16" points="257" swimtime="00:00:39.20" resultid="175810073" heatid="87" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Walkowicz" birthdate="1932-05-18" gender="F" nation="POL" swrid="4877350" athleteid="4877350">
              <RESULTS>
                <RESULT eventid="2" points="14" swimtime="00:01:33.57" resultid="175810070" heatid="16" lane="1" />
                <RESULT eventid="10" points="17" swimtime="00:01:36.90" resultid="175810071" heatid="62" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Mróz" birthdate="1979-06-09" gender="F" nation="POL" swrid="4780617" athleteid="4780617">
              <RESULTS>
                <RESULT eventid="6" points="273" swimtime="00:02:49.94" resultid="175810042" heatid="41" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:21.03" />
                    <SPLIT distance="150" swimtime="00:02:05.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="12" points="230" swimtime="00:01:29.50" resultid="175810041" heatid="69" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Koenig" birthdate="1987-04-21" gender="F" nation="POL" swrid="5464149" athleteid="5464149">
              <RESULTS>
                <RESULT eventid="10" points="47" swimtime="00:01:09.66" resultid="175810054" heatid="61" lane="5" />
                <RESULT eventid="15" points="110" swimtime="00:00:59.55" resultid="175810051" heatid="86" lane="5" />
                <RESULT eventid="17" points="102" swimtime="00:02:13.10" resultid="175810053" heatid="97" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="98" swimtime="00:04:51.65" resultid="175810052" heatid="108" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.94" />
                    <SPLIT distance="100" swimtime="00:02:15.73" />
                    <SPLIT distance="150" swimtime="00:03:31.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Ilnicki" birthdate="1956-03-22" gender="M" nation="POL" swrid="5484406" athleteid="5484406">
              <RESULTS>
                <RESULT eventid="16" points="149" swimtime="00:00:47.01" resultid="175810037" heatid="82" lane="2" />
                <RESULT eventid="18" points="144" swimtime="00:01:45.29" resultid="175810039" heatid="100" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="122" swimtime="00:00:43.76" resultid="175810038" heatid="119" lane="1" />
                <RESULT eventid="30" points="119" swimtime="00:01:39.93" resultid="175810040" heatid="139" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Mrozinski" birthdate="1959-12-28" gender="M" nation="POL" swrid="4877351" athleteid="4877351">
              <RESULTS>
                <RESULT eventid="16" points="329" swimtime="00:00:36.14" resultid="175810055" heatid="87" lane="5" />
                <RESULT eventid="20" points="275" swimtime="00:03:04.71" resultid="175810056" heatid="110" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:01:27.96" />
                    <SPLIT distance="150" swimtime="00:02:15.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jolanta" lastname="Stefanek" birthdate="1960-03-15" gender="F" nation="POL" swrid="4992640" athleteid="4992640">
              <RESULTS>
                <RESULT eventid="15" points="223" swimtime="00:00:47.04" resultid="175810057" heatid="85" lane="4" />
                <RESULT eventid="17" points="198" swimtime="00:01:46.86" resultid="175810059" heatid="98" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="189" swimtime="00:03:54.19" resultid="175810058" heatid="109" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.77" />
                    <SPLIT distance="100" swimtime="00:01:51.58" />
                    <SPLIT distance="150" swimtime="00:02:53.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01203" nation="POL" region="03" clubid="71347" swrid="71347" name="UKS Trójka Puławy" shortname="Trojka Pulawy">
          <ATHLETES>
            <ATHLETE firstname="Witold" lastname="Marciniec" birthdate="1984-03-25" gender="M" nation="POL" swrid="5416820" athleteid="5416820">
              <RESULTS>
                <RESULT eventid="3" points="242" swimtime="00:01:11.88" resultid="175810487" heatid="21" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="265" swimtime="00:05:30.32" resultid="175810488" heatid="46" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:17.58" />
                    <SPLIT distance="150" swimtime="00:01:58.79" />
                    <SPLIT distance="200" swimtime="00:02:40.97" />
                    <SPLIT distance="250" swimtime="00:03:24.08" />
                    <SPLIT distance="300" swimtime="00:04:06.70" />
                    <SPLIT distance="350" swimtime="00:04:47.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Gogacz" birthdate="1976-10-28" gender="M" nation="POL" license="501203700057" swrid="4754646" athleteid="4754646">
              <RESULTS>
                <RESULT eventid="7" points="336" swimtime="00:05:05.18" resultid="175810490" heatid="52" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:14.29" />
                    <SPLIT distance="150" swimtime="00:01:53.42" />
                    <SPLIT distance="200" swimtime="00:02:32.60" />
                    <SPLIT distance="250" swimtime="00:03:10.91" />
                    <SPLIT distance="300" swimtime="00:03:49.50" />
                    <SPLIT distance="350" swimtime="00:04:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="25" points="348" swimtime="00:02:33.76" resultid="175810489" heatid="128" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:13.99" />
                    <SPLIT distance="150" swimtime="00:01:53.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02705" nation="POL" region="05" clubid="86219" swrid="86219" name="TSP Pływak Tomaszów Mazowiecki">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Bucholz" birthdate="1972-01-26" gender="M" nation="POL" swrid="4754642" athleteid="4754642">
              <RESULTS>
                <RESULT eventid="3" points="299" swimtime="00:01:07.00" resultid="175810218" heatid="20" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="289" swimtime="00:02:30.22" resultid="175810216" heatid="42" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="150" swimtime="00:01:52.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="301" swimtime="00:05:16.37" resultid="175810219" heatid="48" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:01:15.63" />
                    <SPLIT distance="150" swimtime="00:01:56.18" />
                    <SPLIT distance="200" swimtime="00:02:37.07" />
                    <SPLIT distance="250" swimtime="00:03:17.22" />
                    <SPLIT distance="300" swimtime="00:03:57.05" />
                    <SPLIT distance="350" swimtime="00:04:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" points="248" swimtime="00:02:54.28" resultid="175810217" heatid="132" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                    <SPLIT distance="100" swimtime="00:01:26.39" />
                    <SPLIT distance="150" swimtime="00:02:16.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00908" nation="POL" region="08" clubid="78661" swrid="78661" name="SP MOTYL przy MOSiR Stalowa Wola" shortname="SP MOTYL MOSiR Stalowa Wola">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Petecka" birthdate="1967-04-17" gender="F" nation="POL" swrid="4992840" athleteid="4992840">
              <RESULTS>
                <RESULT eventid="2" points="249" swimtime="00:00:36.40" resultid="175809966" heatid="9" lane="3" />
                <RESULT eventid="21" points="217" swimtime="00:00:40.57" resultid="175809968" heatid="116" lane="3" />
                <RESULT eventid="27" points="229" swimtime="00:03:18.92" resultid="175809967" heatid="134" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                    <SPLIT distance="100" swimtime="00:01:38.03" />
                    <SPLIT distance="150" swimtime="00:02:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="233" swimtime="00:01:31.75" resultid="175809969" heatid="143" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arkadiusz" lastname="Berwecki" birthdate="1973-01-14" gender="M" nation="POL" license="100908700263" swrid="4791744" athleteid="4791744">
              <RESULTS>
                <RESULT eventid="5" points="482" swimtime="00:02:06.68" resultid="175809962" heatid="39" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="100" swimtime="00:01:01.88" />
                    <SPLIT distance="150" swimtime="00:01:34.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="459" swimtime="00:04:34.96" resultid="175809965" heatid="50" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="150" swimtime="00:01:42.37" />
                    <SPLIT distance="200" swimtime="00:02:17.84" />
                    <SPLIT distance="250" swimtime="00:02:52.89" />
                    <SPLIT distance="300" swimtime="00:03:27.71" />
                    <SPLIT distance="350" swimtime="00:04:02.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" points="443" swimtime="00:01:02.66" resultid="175809963" heatid="125" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="25" points="419" swimtime="00:02:24.61" resultid="175809964" heatid="130" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:10.05" />
                    <SPLIT distance="150" swimtime="00:01:47.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" region="14" clubid="67908" swrid="67908" name="UKS DELFIN Legionowo">
          <ATHLETES>
            <ATHLETE firstname="Joanna" lastname="Żbikowska" birthdate="1996-01-31" gender="F" nation="POL" swrid="4605445" athleteid="4605445">
              <RESULTS>
                <RESULT eventid="15" points="459" swimtime="00:00:37.00" resultid="175810074" heatid="88" lane="1" />
                <RESULT eventid="17" points="458" swimtime="00:01:20.85" resultid="175810076" heatid="101" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="425" swimtime="00:02:58.91" resultid="175810075" heatid="112" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:27.17" />
                    <SPLIT distance="150" swimtime="00:02:13.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="439" swimtime="00:01:14.32" resultid="175810077" heatid="138" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="77480" swrid="77480" name="Warsaw Masters Team">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Giejsztowt" birthdate="1978-06-13" gender="M" nation="POL" swrid="5241012" athleteid="5241012">
              <RESULTS>
                <RESULT eventid="1" points="380" swimtime="00:00:27.81" resultid="175810133" heatid="18" lane="2" />
                <RESULT eventid="3" points="411" swimtime="00:01:00.29" resultid="175810135" heatid="34" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="413" swimtime="00:02:13.35" resultid="175810134" heatid="39" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:01:03.92" />
                    <SPLIT distance="150" swimtime="00:01:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="401" swimtime="00:04:47.65" resultid="175810136" heatid="52" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:07.54" />
                    <SPLIT distance="150" swimtime="00:01:43.23" />
                    <SPLIT distance="200" swimtime="00:02:20.33" />
                    <SPLIT distance="250" swimtime="00:02:57.42" />
                    <SPLIT distance="300" swimtime="00:03:35.19" />
                    <SPLIT distance="350" swimtime="00:04:12.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dymitr" lastname="Bielski" birthdate="1977-08-13" gender="M" nation="POL" swrid="5552366" athleteid="5552366">
              <RESULTS>
                <RESULT eventid="3" points="265" swimtime="00:01:09.80" resultid="175810109" heatid="28" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="295" swimtime="00:02:29.15" resultid="175810107" heatid="42" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:12.08" />
                    <SPLIT distance="150" swimtime="00:01:50.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="276" swimtime="00:05:25.84" resultid="175810110" heatid="48" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:15.06" />
                    <SPLIT distance="150" swimtime="00:01:55.71" />
                    <SPLIT distance="200" swimtime="00:03:19.27" />
                    <SPLIT distance="250" swimtime="00:04:01.80" />
                    <SPLIT distance="300" swimtime="00:04:44.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="320" swimtime="00:02:55.53" resultid="175810108" heatid="110" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:01:24.41" />
                    <SPLIT distance="150" swimtime="00:02:09.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ostrowski" birthdate="1977-05-14" gender="M" nation="POL" license="504214700091" swrid="5506635" athleteid="5506635">
              <RESULTS>
                <RESULT eventid="3" points="434" swimtime="00:00:59.21" resultid="175810117" heatid="33" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="340" swimtime="00:05:03.90" resultid="175810118" heatid="48" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:50.04" />
                    <SPLIT distance="200" swimtime="00:02:27.96" />
                    <SPLIT distance="250" swimtime="00:03:06.71" />
                    <SPLIT distance="300" swimtime="00:03:45.57" />
                    <SPLIT distance="350" swimtime="00:04:22.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="488" swimtime="00:00:31.68" resultid="175810115" heatid="89" lane="1" />
                <RESULT eventid="20" points="352" swimtime="00:02:50.17" resultid="175810116" heatid="105" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:21.41" />
                    <SPLIT distance="150" swimtime="00:02:05.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafal" lastname="Skoskiewicz" birthdate="1966-05-05" gender="M" nation="POL" license="504214700002" swrid="4183802" athleteid="4183802">
              <RESULTS>
                <RESULT eventid="7" points="410" swimtime="00:04:45.55" resultid="175810132" heatid="52" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="100" swimtime="00:01:08.10" />
                    <SPLIT distance="150" swimtime="00:01:44.27" />
                    <SPLIT distance="200" swimtime="00:02:21.15" />
                    <SPLIT distance="250" swimtime="00:02:58.38" />
                    <SPLIT distance="300" swimtime="00:03:35.16" />
                    <SPLIT distance="350" swimtime="00:04:10.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11" points="366" swimtime="00:01:07.55" resultid="175810129" heatid="70" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" points="377" swimtime="00:02:31.65" resultid="175810130" heatid="136" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                    <SPLIT distance="150" swimtime="00:01:56.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="376" swimtime="00:01:08.24" resultid="175810131" heatid="142" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pawel" lastname="Rogosz" birthdate="1976-04-28" gender="M" nation="POL" license="504214700003" swrid="4270348" athleteid="4270348">
              <RESULTS>
                <RESULT eventid="11" points="259" swimtime="00:01:15.80" resultid="175810111" heatid="67" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" points="364" swimtime="00:01:17.40" resultid="175810113" heatid="96" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="377" swimtime="00:02:46.29" resultid="175810112" heatid="105" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:21.24" />
                    <SPLIT distance="150" swimtime="00:02:04.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="25" points="293" swimtime="00:02:42.92" resultid="175810114" heatid="128" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:20.14" />
                    <SPLIT distance="150" swimtime="00:02:01.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miroslaw" lastname="Warchol" birthdate="1953-08-30" gender="M" nation="POL" swrid="4222718" athleteid="4222718">
              <RESULTS>
                <RESULT eventid="11" points="218" swimtime="00:01:20.30" resultid="175810119" heatid="67" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="236" swimtime="00:02:50.80" resultid="175810120" heatid="73" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:22.64" />
                    <SPLIT distance="150" swimtime="00:02:06.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Bielecka" birthdate="1988-04-07" gender="F" nation="POL" swrid="5582449" athleteid="5582449">
              <RESULTS>
                <RESULT eventid="15" points="384" swimtime="00:00:39.27" resultid="175810121" heatid="88" lane="6" />
                <RESULT eventid="21" points="333" swimtime="00:00:35.17" resultid="175810123" heatid="113" lane="1" />
                <RESULT eventid="26" points="271" swimtime="00:03:04.70" resultid="175810124" heatid="129" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:15.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="27" points="369" swimtime="00:02:49.88" resultid="175810122" heatid="131" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:19.48" />
                    <SPLIT distance="150" swimtime="00:02:08.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Porada" birthdate="1983-06-10" gender="M" nation="POL" swrid="5506638" athleteid="5506638">
              <RESULTS>
                <RESULT eventid="16" points="437" swimtime="00:00:32.86" resultid="175810125" heatid="84" lane="3" />
                <RESULT eventid="20" points="406" swimtime="00:02:42.27" resultid="175810126" heatid="105" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                    <SPLIT distance="150" swimtime="00:01:59.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="402" swimtime="00:00:29.45" resultid="175810127" heatid="120" lane="2" />
                <RESULT eventid="25" points="349" swimtime="00:02:33.73" resultid="175810128" heatid="128" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="150" swimtime="00:01:51.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00706" nation="POL" region="06" clubid="74345" swrid="74345" name="UKS SP 8 Chrzanów">
          <ATHLETES>
            <ATHLETE firstname="Alfred" lastname="Zabrzański" birthdate="1954-05-12" gender="M" nation="POL" swrid="4477631" athleteid="4477631">
              <RESULTS>
                <RESULT eventid="1" points="222" swimtime="00:00:33.28" resultid="175810139" heatid="7" lane="4" />
                <RESULT eventid="3" points="208" swimtime="00:01:15.58" resultid="175810141" heatid="25" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="180" swimtime="00:02:55.93" resultid="175810140" heatid="43" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:24.13" />
                    <SPLIT distance="150" swimtime="00:02:10.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="132" swimtime="00:00:43.62" resultid="175810142" heatid="57" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00111" nation="POL" region="11" clubid="65944" swrid="65944" name="UKS TRÓJKA Częstochowa">
          <ATHLETES>
            <ATHLETE firstname="Wiktoria" lastname="Musik" birthdate="1997-08-04" gender="F" nation="POL" license="100111600053" swrid="4602697" athleteid="4602697">
              <RESULTS>
                <RESULT eventid="2" points="585" swimtime="00:00:27.41" resultid="175810465" heatid="15" lane="3" />
                <RESULT eventid="4" points="584" swimtime="00:01:00.11" resultid="175810467" heatid="23" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" points="538" swimtime="00:02:15.59" resultid="175810466" heatid="37" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="100" swimtime="00:01:04.32" />
                    <SPLIT distance="150" swimtime="00:01:40.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="547" swimtime="00:01:09.09" resultid="175810468" heatid="146" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Warwas" birthdate="1995-07-13" gender="M" nation="POL" swrid="4266133" athleteid="4266133">
              <RESULTS>
                <RESULT eventid="1" points="497" swimtime="00:00:25.45" resultid="175810477" heatid="13" lane="2" />
                <RESULT eventid="9" points="369" swimtime="00:00:30.97" resultid="175810480" heatid="59" lane="2" />
                <RESULT eventid="22" points="446" swimtime="00:00:28.45" resultid="175810479" heatid="122" lane="4" />
                <RESULT eventid="24" points="330" swimtime="00:01:09.09" resultid="175810478" heatid="127" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Gajda" birthdate="1995-04-24" gender="M" nation="POL" license="100111700062" swrid="4762175" athleteid="4762175">
              <RESULTS>
                <RESULT eventid="1" points="543" swimtime="00:00:24.71" resultid="175810481" heatid="8" lane="4" />
                <RESULT eventid="3" points="521" swimtime="00:00:55.71" resultid="175810484" heatid="30" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="527" swimtime="00:00:26.92" resultid="175810483" heatid="117" lane="4" />
                <RESULT eventid="24" points="512" swimtime="00:00:59.69" resultid="175810482" heatid="125" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kurek" birthdate="1994-07-11" gender="M" nation="POL" license="100111700097" swrid="5502059" athleteid="5502059">
              <RESULTS>
                <RESULT eventid="3" points="387" swimtime="00:01:01.50" resultid="175810471" heatid="34" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="347" swimtime="00:00:35.48" resultid="175810469" heatid="87" lane="3" />
                <RESULT eventid="28" points="309" swimtime="00:02:42.03" resultid="175810470" heatid="136" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:14.52" />
                    <SPLIT distance="150" swimtime="00:02:01.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="343" swimtime="00:01:10.36" resultid="175810472" heatid="147" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sonia" lastname="Nowak" birthdate="1996-05-23" gender="F" nation="POL" license="100111600092" swrid="4289072" athleteid="4289072">
              <RESULTS>
                <RESULT eventid="6" points="457" swimtime="00:02:23.11" resultid="175810473" heatid="37" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:07.33" />
                    <SPLIT distance="150" swimtime="00:01:44.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8" points="453" swimtime="00:05:04.42" resultid="175810476" heatid="53" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                    <SPLIT distance="150" swimtime="00:01:53.90" />
                    <SPLIT distance="200" swimtime="00:02:32.65" />
                    <SPLIT distance="250" swimtime="00:03:11.30" />
                    <SPLIT distance="300" swimtime="00:03:49.64" />
                    <SPLIT distance="350" swimtime="00:04:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" points="405" swimtime="00:01:13.78" resultid="175810474" heatid="123" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="26" points="410" swimtime="00:02:40.93" resultid="175810475" heatid="129" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:16.60" />
                    <SPLIT distance="150" swimtime="00:01:58.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="31" points="535" swimtime="00:01:48.22" resultid="175810485" heatid="150" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.53" />
                    <SPLIT distance="100" swimtime="00:00:58.22" />
                    <SPLIT distance="150" swimtime="00:01:23.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4602697" number="1" />
                    <RELAYPOSITION athleteid="4289072" number="2" />
                    <RELAYPOSITION athleteid="4266133" number="3" />
                    <RELAYPOSITION athleteid="4762175" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="445" swimtime="00:02:05.92" resultid="175810486" heatid="152" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                    <SPLIT distance="150" swimtime="00:01:34.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4602697" number="1" />
                    <RELAYPOSITION athleteid="5502059" number="2" />
                    <RELAYPOSITION athleteid="4762175" number="3" />
                    <RELAYPOSITION athleteid="4289072" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="08001" nation="POL" region="01" clubid="93972" swrid="93972" name="Sport Active">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Mroczko" birthdate="1978-01-30" gender="M" nation="POL" swrid="5626922" athleteid="5626922">
              <RESULTS>
                <RESULT eventid="1" points="169" swimtime="00:00:36.42" resultid="175809846" heatid="3" lane="6" />
                <RESULT eventid="3" points="157" swimtime="00:01:23.00" resultid="175809848" heatid="21" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="151" swimtime="00:03:06.26" resultid="175809847" heatid="36" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                    <SPLIT distance="100" swimtime="00:01:28.57" />
                    <SPLIT distance="150" swimtime="00:02:17.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="146" swimtime="00:06:42.77" resultid="175809849" heatid="46" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                    <SPLIT distance="100" swimtime="00:01:32.09" />
                    <SPLIT distance="150" swimtime="00:02:23.64" />
                    <SPLIT distance="200" swimtime="00:03:15.77" />
                    <SPLIT distance="250" swimtime="00:04:08.95" />
                    <SPLIT distance="300" swimtime="00:05:02.24" />
                    <SPLIT distance="350" swimtime="00:05:54.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Cygal" birthdate="1980-09-10" gender="M" nation="POL" swrid="5626900" athleteid="5626900">
              <RESULTS>
                <RESULT eventid="1" points="150" swimtime="00:00:37.89" resultid="175809852" heatid="3" lane="2" />
                <RESULT eventid="7" points="98" swimtime="00:07:39.59" resultid="175809855" heatid="46" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.78" />
                    <SPLIT distance="100" swimtime="00:01:40.87" />
                    <SPLIT distance="150" swimtime="00:02:37.93" />
                    <SPLIT distance="200" swimtime="00:03:37.98" />
                    <SPLIT distance="250" swimtime="00:04:40.26" />
                    <SPLIT distance="300" swimtime="00:05:43.32" />
                    <SPLIT distance="350" swimtime="00:06:43.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" points="155" swimtime="00:01:42.90" resultid="175809854" heatid="93" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="150" swimtime="00:03:46.01" resultid="175809853" heatid="103" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                    <SPLIT distance="100" swimtime="00:01:46.70" />
                    <SPLIT distance="150" swimtime="00:02:48.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Cygal" birthdate="1981-09-17" gender="F" nation="POL" swrid="5626899" athleteid="5626899">
              <RESULTS>
                <RESULT eventid="15" points="121" swimtime="00:00:57.71" resultid="175809840" heatid="77" lane="4" />
                <RESULT eventid="17" points="101" swimtime="00:02:13.63" resultid="175809842" heatid="91" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="103" swimtime="00:04:46.32" resultid="175809841" heatid="102" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.99" />
                    <SPLIT distance="100" swimtime="00:02:17.63" />
                    <SPLIT distance="150" swimtime="00:03:33.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Wiatrowska" birthdate="1977-08-28" gender="F" nation="POL" swrid="5626944" athleteid="5626944">
              <RESULTS>
                <RESULT eventid="15" points="83" swimtime="00:01:05.41" resultid="175809843" heatid="78" lane="2" />
                <RESULT eventid="17" points="90" swimtime="00:02:18.67" resultid="175809845" heatid="92" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="76" swimtime="00:05:17.10" resultid="175809844" heatid="102" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.76" />
                    <SPLIT distance="100" swimtime="00:02:24.72" />
                    <SPLIT distance="150" swimtime="00:03:51.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="31" points="99" swimtime="00:03:09.55" resultid="175809850" heatid="148" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.50" />
                    <SPLIT distance="100" swimtime="00:01:55.21" />
                    <SPLIT distance="150" swimtime="00:02:32.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5626944" number="1" />
                    <RELAYPOSITION athleteid="5626899" number="2" />
                    <RELAYPOSITION athleteid="5626900" number="3" />
                    <RELAYPOSITION athleteid="5626922" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="84" swimtime="00:03:38.90" resultid="175809851" heatid="152" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.68" />
                    <SPLIT distance="100" swimtime="00:02:13.59" />
                    <SPLIT distance="150" swimtime="00:03:01.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5626944" number="1" />
                    <RELAYPOSITION athleteid="5626899" number="2" />
                    <RELAYPOSITION athleteid="5626900" number="3" />
                    <RELAYPOSITION athleteid="5626922" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="NATION" code="CZE" nation="CZE" clubid="94" swrid="94" name="Czech Republic">
          <ATHLETES>
            <ATHLETE firstname="Vaclav" lastname="Valtr" birthdate="1956-07-10" gender="M" nation="CZE" swrid="4182881" athleteid="4182881">
              <RESULTS>
                <RESULT eventid="3" points="252" swimtime="00:01:10.98" resultid="175810345" heatid="28" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11" points="217" swimtime="00:01:20.34" resultid="175810343" heatid="67" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="203" swimtime="00:03:24.14" resultid="175810344" heatid="107" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="100" swimtime="00:01:39.67" />
                    <SPLIT distance="150" swimtime="00:02:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="234" swimtime="00:01:19.96" resultid="175810346" heatid="144" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dana" lastname="Benova" birthdate="1956-01-26" gender="F" nation="CZE" swrid="4223032" athleteid="4223032">
              <RESULTS>
                <RESULT eventid="6" points="65" swimtime="00:04:33.75" resultid="175810339" heatid="41" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.58" />
                    <SPLIT distance="100" swimtime="00:02:09.74" />
                    <SPLIT distance="150" swimtime="00:03:22.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8" points="66" swimtime="00:09:36.59" resultid="175810342" heatid="49" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.77" />
                    <SPLIT distance="100" swimtime="00:02:15.07" />
                    <SPLIT distance="150" swimtime="00:03:30.19" />
                    <SPLIT distance="200" swimtime="00:04:45.66" />
                    <SPLIT distance="250" swimtime="00:05:59.28" />
                    <SPLIT distance="300" swimtime="00:07:13.18" />
                    <SPLIT distance="350" swimtime="00:08:27.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="17" points="72" swimtime="00:02:29.35" resultid="175810341" heatid="97" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="83" swimtime="00:05:07.75" resultid="175810340" heatid="111" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.52" />
                    <SPLIT distance="100" swimtime="00:02:35.96" />
                    <SPLIT distance="150" swimtime="00:03:55.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00601" nation="POL" region="01" clubid="65965" swrid="65965" name="WKS ŚLĄSK Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Rother" birthdate="1968-05-21" gender="M" nation="POL" swrid="4351633" athleteid="4351633">
              <RESULTS>
                <RESULT eventid="9" points="358" swimtime="00:00:31.29" resultid="175810080" heatid="59" lane="5" />
                <RESULT eventid="11" points="349" swimtime="00:01:08.59" resultid="175810078" heatid="70" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="341" swimtime="00:02:31.15" resultid="175810079" heatid="73" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:14.87" />
                    <SPLIT distance="150" swimtime="00:01:52.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01012" nation="POL" region="12" clubid="86431" swrid="86431" name="MOSiR Ostrowiec Świętokrzyski" shortname="MOSiR Ostrowiec">
          <ATHLETES>
            <ATHLETE firstname="Jósef" lastname="Rózalski" birthdate="1945-03-28" gender="M" nation="POL" swrid="4216999" athleteid="4216999">
              <RESULTS>
                <RESULT eventid="16" points="66" swimtime="00:01:01.55" resultid="175810464" heatid="90" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="NATION" code="POL" nation="POL" clubid="291" swrid="291" name="Poland">
          <ATHLETES>
            <ATHLETE firstname="Marta" lastname="Czarnecka" birthdate="2002-08-27" gender="F" nation="POL" swrid="5175088" athleteid="5175088">
              <RESULTS>
                <RESULT eventid="2" points="346" swimtime="00:00:32.64" resultid="175810244" heatid="4" lane="1" />
                <RESULT eventid="15" points="386" swimtime="00:00:39.22" resultid="175810243" heatid="80" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Rudzki" birthdate="1992-06-21" gender="M" nation="POL" swrid="4250678" athleteid="4250678">
              <RESULTS>
                <RESULT eventid="1" points="423" swimtime="00:00:26.85" resultid="175810555" heatid="8" lane="5" />
                <RESULT eventid="3" points="448" swimtime="00:00:58.58" resultid="175810557" heatid="30" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" points="413" swimtime="00:02:27.12" resultid="175810556" heatid="136" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                    <SPLIT distance="100" swimtime="00:01:06.84" />
                    <SPLIT distance="150" swimtime="00:01:50.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="426" swimtime="00:01:05.47" resultid="175810558" heatid="142" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Źródlak" birthdate="1997-10-31" gender="M" nation="POL" swrid="4288152" athleteid="4288152">
              <RESULTS>
                <RESULT eventid="1" points="302" swimtime="00:00:30.02" resultid="175810547" heatid="7" lane="1" />
                <RESULT eventid="9" points="220" swimtime="00:00:36.80" resultid="175810550" heatid="55" lane="6" />
                <RESULT eventid="16" points="214" swimtime="00:00:41.71" resultid="175810548" heatid="83" lane="6" />
                <RESULT eventid="18" points="237" swimtime="00:01:29.22" resultid="175810549" heatid="94" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Bart" birthdate="1997-10-10" gender="F" nation="POL" swrid="4289388" athleteid="4289388">
              <RESULTS>
                <RESULT eventid="2" points="513" swimtime="00:00:28.63" resultid="175810565" heatid="5" lane="6" />
                <RESULT eventid="4" points="481" swimtime="00:01:04.12" resultid="175810568" heatid="23" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" points="529" swimtime="00:02:16.33" resultid="175810566" heatid="45" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                    <SPLIT distance="150" swimtime="00:01:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" points="447" swimtime="00:00:31.87" resultid="175810567" heatid="118" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Gajdowski" birthdate="1988-10-10" gender="M" nation="POL" swrid="4369675" athleteid="4369675">
              <RESULTS>
                <RESULT eventid="1" points="380" swimtime="00:00:27.81" resultid="175810261" heatid="12" lane="4" />
                <RESULT eventid="16" points="311" swimtime="00:00:36.82" resultid="175810262" heatid="84" lane="1" />
                <RESULT eventid="18" points="328" swimtime="00:01:20.14" resultid="175810263" heatid="96" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="314" swimtime="00:01:12.50" resultid="175810264" heatid="147" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Kutyło" birthdate="1999-02-13" gender="F" nation="POL" swrid="4496783" athleteid="4496783">
              <RESULTS>
                <RESULT eventid="2" points="368" swimtime="00:00:31.98" resultid="175810347" heatid="9" lane="4" />
                <RESULT eventid="6" points="281" swimtime="00:02:48.40" resultid="175810348" heatid="38" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                    <SPLIT distance="100" swimtime="00:01:22.08" />
                    <SPLIT distance="150" swimtime="00:02:06.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" points="297" swimtime="00:00:36.54" resultid="175810349" heatid="118" lane="1" />
                <RESULT eventid="29" points="300" swimtime="00:01:24.35" resultid="175810350" heatid="137" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Apolonia" lastname="Popławska" birthdate="2002-06-01" gender="F" nation="POL" license="100515600277" swrid="4946114" athleteid="4946114">
              <RESULTS>
                <RESULT eventid="2" points="485" swimtime="00:00:29.17" resultid="175810522" heatid="15" lane="2" />
                <RESULT eventid="15" points="503" swimtime="00:00:35.90" resultid="175810523" heatid="88" lane="3" />
                <RESULT eventid="21" points="463" swimtime="00:00:31.51" resultid="175810524" heatid="113" lane="4" />
                <RESULT eventid="29" points="496" swimtime="00:01:11.38" resultid="175810525" heatid="146" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Poppe" birthdate="2003-08-28" gender="F" nation="POL" swrid="5062765" athleteid="5062765">
              <RESULTS>
                <RESULT eventid="2" points="419" swimtime="00:00:30.63" resultid="175810331" heatid="4" lane="3" />
                <RESULT eventid="19" points="347" swimtime="00:03:11.42" resultid="175810332" heatid="112" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:28.71" />
                    <SPLIT distance="150" swimtime="00:02:18.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ryszard" lastname="Zając" birthdate="1984-07-29" gender="M" nation="POL" swrid="5468089" athleteid="5468089">
              <RESULTS>
                <RESULT eventid="1" points="180" swimtime="00:00:35.65" resultid="175810290" heatid="11" lane="4" />
                <RESULT eventid="3" points="179" swimtime="00:01:19.47" resultid="175810292" heatid="25" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="161" swimtime="00:00:45.86" resultid="175810291" heatid="90" lane="1" />
                <RESULT eventid="30" points="128" swimtime="00:01:37.64" resultid="175810293" heatid="141" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Jania" birthdate="1988-01-01" gender="M" nation="POL" swrid="5484407" athleteid="5484407">
              <RESULTS>
                <RESULT eventid="1" points="190" swimtime="00:00:35.03" resultid="175810294" heatid="19" lane="2" />
                <RESULT eventid="16" points="189" swimtime="00:00:43.45" resultid="175810295" heatid="79" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Jasik" birthdate="1984-01-01" gender="F" nation="POL" swrid="5484408" athleteid="5484408">
              <RESULTS>
                <RESULT eventid="2" points="261" swimtime="00:00:35.86" resultid="175810286" heatid="5" lane="4" />
                <RESULT eventid="4" points="230" swimtime="00:01:21.90" resultid="175810288" heatid="22" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" points="233" swimtime="00:02:59.14" resultid="175810287" heatid="45" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                    <SPLIT distance="100" swimtime="00:01:21.86" />
                    <SPLIT distance="150" swimtime="00:02:09.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8" points="224" swimtime="00:06:25.14" resultid="175810289" heatid="49" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                    <SPLIT distance="100" swimtime="00:01:25.29" />
                    <SPLIT distance="150" swimtime="00:02:13.60" />
                    <SPLIT distance="200" swimtime="00:03:03.74" />
                    <SPLIT distance="250" swimtime="00:03:54.28" />
                    <SPLIT distance="300" swimtime="00:04:45.29" />
                    <SPLIT distance="350" swimtime="00:05:37.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Piórkowski" birthdate="1965-07-28" gender="M" nation="POL" license="510414700072" swrid="5506637" athleteid="5506637">
              <RESULTS>
                <RESULT eventid="1" points="140" swimtime="00:00:38.79" resultid="175810306" heatid="19" lane="5" />
                <RESULT eventid="3" points="143" swimtime="00:01:25.61" resultid="175810308" heatid="29" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="128" swimtime="00:03:16.89" resultid="175810307" heatid="44" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                    <SPLIT distance="100" swimtime="00:01:33.25" />
                    <SPLIT distance="150" swimtime="00:02:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="98" swimtime="00:00:48.19" resultid="175810309" heatid="56" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Sarna" birthdate="1975-10-31" gender="M" nation="POL" swrid="5540150" athleteid="5540150">
              <RESULTS>
                <RESULT eventid="1" points="397" swimtime="00:00:27.41" resultid="175810573" heatid="12" lane="1" />
                <RESULT eventid="3" points="413" swimtime="00:01:00.19" resultid="175810575" heatid="33" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="411" swimtime="00:02:13.56" resultid="175810574" heatid="39" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                    <SPLIT distance="100" swimtime="00:01:02.22" />
                    <SPLIT distance="150" swimtime="00:01:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="345" swimtime="00:01:10.25" resultid="175810576" heatid="147" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Batóg" birthdate="1972-03-11" gender="F" nation="POL" swrid="5626895" athleteid="5626895">
              <RESULTS>
                <RESULT eventid="2" points="293" swimtime="00:00:34.50" resultid="175810318" heatid="5" lane="2" />
                <RESULT eventid="21" points="219" swimtime="00:00:40.44" resultid="175810320" heatid="118" lane="4" />
                <RESULT eventid="23" points="215" swimtime="00:01:31.10" resultid="175810319" heatid="123" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="264" swimtime="00:01:27.99" resultid="175810321" heatid="137" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Broniszewski" birthdate="1980-09-29" gender="M" nation="POL" swrid="5626896" athleteid="5626896">
              <RESULTS>
                <RESULT eventid="1" points="231" swimtime="00:00:32.85" resultid="175810539" heatid="7" lane="6" />
                <RESULT eventid="3" points="216" swimtime="00:01:14.62" resultid="175810541" heatid="25" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="231" swimtime="00:00:40.62" resultid="175810540" heatid="83" lane="2" />
                <RESULT eventid="18" points="239" swimtime="00:01:29.00" resultid="175810542" heatid="99" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Bukowski" birthdate="1981-01-01" gender="M" nation="POL" swrid="5626897" athleteid="5626897">
              <RESULTS>
                <RESULT eventid="1" points="343" swimtime="00:00:28.79" resultid="175810300" heatid="12" lane="2" />
                <RESULT eventid="20" points="270" swimtime="00:03:05.77" resultid="175810301" heatid="104" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:29.25" />
                    <SPLIT distance="150" swimtime="00:02:17.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="324" swimtime="00:00:31.65" resultid="175810302" heatid="120" lane="3" />
                <RESULT eventid="30" points="272" swimtime="00:01:15.98" resultid="175810303" heatid="144" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Faff" birthdate="1963-01-01" gender="M" nation="POL" swrid="5626904" athleteid="5626904">
              <RESULTS>
                <RESULT eventid="1" points="305" swimtime="00:00:29.94" resultid="175810577" heatid="17" lane="3" />
                <RESULT eventid="3" points="298" swimtime="00:01:07.12" resultid="175810580" heatid="20" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="251" swimtime="00:02:37.52" resultid="175810578" heatid="35" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:13.51" />
                    <SPLIT distance="150" swimtime="00:01:56.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="266" swimtime="00:00:33.79" resultid="175810579" heatid="120" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Kapera" birthdate="1967-06-20" gender="M" nation="POL" swrid="5626908" athleteid="5626908">
              <RESULTS>
                <RESULT eventid="1" points="168" swimtime="00:00:36.53" resultid="175810569" heatid="3" lane="5" />
                <RESULT eventid="3" points="153" swimtime="00:01:23.82" resultid="175810572" heatid="31" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="142" swimtime="00:03:10.38" resultid="175810570" heatid="40" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                    <SPLIT distance="100" swimtime="00:01:30.42" />
                    <SPLIT distance="150" swimtime="00:02:21.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="118" swimtime="00:00:44.32" resultid="175810571" heatid="121" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Ludynia" birthdate="1979-10-23" gender="M" nation="POL" swrid="5626916" athleteid="5626916">
              <RESULTS>
                <RESULT eventid="1" points="285" swimtime="00:00:30.62" resultid="175810563" heatid="17" lane="6" />
                <RESULT eventid="28" points="213" swimtime="00:03:03.42" resultid="175810564" heatid="132" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                    <SPLIT distance="100" swimtime="00:01:27.02" />
                    <SPLIT distance="150" swimtime="00:02:18.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Marszałek" birthdate="1954-10-24" gender="M" nation="POL" swrid="5626919" athleteid="5626919">
              <RESULTS>
                <RESULT eventid="1" points="106" swimtime="00:00:42.48" resultid="175810518" heatid="19" lane="6" />
                <RESULT eventid="5" points="97" swimtime="00:03:36.07" resultid="175810519" heatid="44" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.15" />
                    <SPLIT distance="100" swimtime="00:01:45.64" />
                    <SPLIT distance="150" swimtime="00:02:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="103" swimtime="00:07:31.74" resultid="175810521" heatid="54" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.88" />
                    <SPLIT distance="100" swimtime="00:01:47.73" />
                    <SPLIT distance="150" swimtime="00:02:45.76" />
                    <SPLIT distance="200" swimtime="00:03:40.81" />
                    <SPLIT distance="250" swimtime="00:04:39.67" />
                    <SPLIT distance="300" swimtime="00:05:35.64" />
                    <SPLIT distance="350" swimtime="00:06:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="67" swimtime="00:00:53.48" resultid="175810520" heatid="115" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Michalczuk" birthdate="1970-03-05" gender="M" nation="POL" swrid="5626920" athleteid="5626920">
              <RESULTS>
                <RESULT eventid="1" points="216" swimtime="00:00:33.58" resultid="175810322" heatid="7" lane="3" />
                <RESULT eventid="3" points="198" swimtime="00:01:16.88" resultid="175810323" heatid="25" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="126" swimtime="00:00:44.27" resultid="175810324" heatid="57" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Miler" birthdate="2002-11-13" gender="M" nation="POL" swrid="5626921" athleteid="5626921">
              <RESULTS>
                <RESULT eventid="1" points="263" swimtime="00:00:31.43" resultid="175810333" heatid="6" lane="2" />
                <RESULT eventid="3" points="254" swimtime="00:01:10.78" resultid="175810336" heatid="28" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="224" swimtime="00:02:43.41" resultid="175810334" heatid="35" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:17.80" />
                    <SPLIT distance="150" swimtime="00:02:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="270" swimtime="00:00:33.65" resultid="175810335" heatid="114" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Niedźwiadek" birthdate="1993-10-18" gender="M" nation="POL" swrid="5626925" athleteid="5626925">
              <RESULTS>
                <RESULT eventid="1" points="344" swimtime="00:00:28.77" resultid="175810543" heatid="18" lane="4" />
                <RESULT eventid="3" points="366" swimtime="00:01:02.66" resultid="175810545" heatid="34" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="357" swimtime="00:02:20.03" resultid="175810544" heatid="39" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="100" swimtime="00:01:06.89" />
                    <SPLIT distance="150" swimtime="00:01:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="404" swimtime="00:04:46.88" resultid="175810546" heatid="52" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:05.75" />
                    <SPLIT distance="150" swimtime="00:01:41.46" />
                    <SPLIT distance="200" swimtime="00:02:17.91" />
                    <SPLIT distance="250" swimtime="00:02:54.77" />
                    <SPLIT distance="300" swimtime="00:03:31.91" />
                    <SPLIT distance="350" swimtime="00:04:09.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iwona" lastname="Nowak" birthdate="1988-01-01" gender="F" nation="POL" swrid="5626926" athleteid="5626926">
              <RESULTS>
                <RESULT eventid="2" points="255" swimtime="00:00:36.13" resultid="175810296" heatid="5" lane="1" />
                <RESULT eventid="10" points="186" swimtime="00:00:44.21" resultid="175810299" heatid="58" lane="1" />
                <RESULT eventid="12" points="186" swimtime="00:01:36.15" resultid="175810297" heatid="65" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="212" swimtime="00:01:34.68" resultid="175810298" heatid="143" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sabina" lastname="Pakosz" birthdate="1981-07-15" gender="F" nation="POL" swrid="5626928" athleteid="5626928">
              <RESULTS>
                <RESULT eventid="2" points="267" swimtime="00:00:35.58" resultid="175810249" heatid="5" lane="5" />
                <RESULT eventid="4" points="255" swimtime="00:01:19.19" resultid="175810250" heatid="22" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Glib" lastname="Pronskikh" birthdate="1991-01-01" gender="M" nation="POL" swrid="5626931" athleteid="5626931">
              <RESULTS>
                <RESULT eventid="1" points="258" swimtime="00:00:31.65" resultid="175810268" heatid="11" lane="1" />
                <RESULT eventid="3" points="185" swimtime="00:01:18.58" resultid="175810270" heatid="24" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="199" swimtime="00:02:50.08" resultid="175810269" heatid="43" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:01:16.88" />
                    <SPLIT distance="150" swimtime="00:02:04.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Szymański" birthdate="1978-01-02" gender="M" nation="POL" swrid="5626939" athleteid="5626939">
              <RESULTS>
                <RESULT eventid="1" points="285" swimtime="00:00:30.62" resultid="175810526" heatid="18" lane="6" />
                <RESULT eventid="3" points="326" swimtime="00:01:05.10" resultid="175810527" heatid="20" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="252" swimtime="00:00:35.15" resultid="175810528" heatid="57" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Wańha" birthdate="1983-04-19" gender="M" nation="POL" swrid="5626942" athleteid="5626942">
              <RESULTS>
                <RESULT eventid="1" points="325" swimtime="00:00:29.30" resultid="175810533" heatid="17" lane="5" />
                <RESULT eventid="3" points="305" swimtime="00:01:06.61" resultid="175810534" heatid="20" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Wciórka" birthdate="1982-06-10" gender="M" nation="POL" swrid="5626943" athleteid="5626943">
              <RESULTS>
                <RESULT eventid="1" points="363" swimtime="00:00:28.26" resultid="175810251" heatid="12" lane="5" />
                <RESULT eventid="9" points="302" swimtime="00:00:33.10" resultid="175810254" heatid="55" lane="2" />
                <RESULT eventid="11" points="231" swimtime="00:01:18.72" resultid="175810252" heatid="70" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="236" swimtime="00:02:50.75" resultid="175810253" heatid="73" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                    <SPLIT distance="100" swimtime="00:01:22.30" />
                    <SPLIT distance="150" swimtime="00:02:07.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Wiciński" birthdate="1987-04-12" gender="M" nation="POL" swrid="5626945" athleteid="5626945">
              <RESULTS>
                <RESULT eventid="1" points="314" swimtime="00:00:29.64" resultid="175810240" heatid="17" lane="1" />
                <RESULT eventid="22" points="262" swimtime="00:00:33.95" resultid="175810241" heatid="119" lane="3" />
                <RESULT eventid="24" points="221" swimtime="00:01:19.02" resultid="175810239" heatid="124" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="275" swimtime="00:01:15.71" resultid="175810242" heatid="144" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Barnasiuk" birthdate="1992-02-04" gender="M" nation="POL" swrid="4273597" athleteid="4273597">
              <RESULTS>
                <RESULT eventid="3" points="440" swimtime="00:00:58.94" resultid="175810537" heatid="33" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="465" swimtime="00:00:32.20" resultid="175810535" heatid="89" lane="5" />
                <RESULT eventid="28" points="447" swimtime="00:02:23.33" resultid="175810536" heatid="136" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                    <SPLIT distance="100" swimtime="00:01:08.21" />
                    <SPLIT distance="150" swimtime="00:01:49.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="423" swimtime="00:01:05.63" resultid="175810538" heatid="142" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Lippa" birthdate="1946-02-02" gender="F" nation="POL" swrid="5484413" athleteid="5484413">
              <RESULTS>
                <RESULT eventid="4" points="10" swimtime="00:03:48.77" resultid="175810504" heatid="26" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" points="18" swimtime="00:07:00.85" resultid="175810502" heatid="41" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.18" />
                    <SPLIT distance="100" swimtime="00:03:24.33" />
                    <SPLIT distance="150" swimtime="00:05:15.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8" points="23" swimtime="00:13:38.27" resultid="175810505" heatid="51" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.35" />
                    <SPLIT distance="100" swimtime="00:03:12.89" />
                    <SPLIT distance="150" swimtime="00:04:59.39" />
                    <SPLIT distance="200" swimtime="00:06:43.20" />
                    <SPLIT distance="250" swimtime="00:08:27.03" />
                    <SPLIT distance="300" swimtime="00:10:10.22" />
                    <SPLIT distance="350" swimtime="00:11:56.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="23" swimtime="00:07:48.39" resultid="175810503" heatid="111" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:48.88" />
                    <SPLIT distance="100" swimtime="00:03:51.09" />
                    <SPLIT distance="150" swimtime="00:05:50.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kędzior" birthdate="1973-12-08" gender="M" nation="POL" swrid="5626909" athleteid="5626909">
              <RESULTS>
                <RESULT eventid="3" points="215" swimtime="00:01:14.78" resultid="175810237" heatid="24" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="197" swimtime="00:06:04.24" resultid="175810238" heatid="48" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:23.61" />
                    <SPLIT distance="150" swimtime="00:02:07.28" />
                    <SPLIT distance="200" swimtime="00:02:53.77" />
                    <SPLIT distance="250" swimtime="00:03:40.79" />
                    <SPLIT distance="300" swimtime="00:04:29.74" />
                    <SPLIT distance="350" swimtime="00:05:17.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11" points="147" swimtime="00:01:31.50" resultid="175810235" heatid="64" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" points="160" swimtime="00:03:21.65" resultid="175810236" heatid="132" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                    <SPLIT distance="100" swimtime="00:01:31.89" />
                    <SPLIT distance="150" swimtime="00:02:37.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Kęsik" birthdate="1979-09-21" gender="M" nation="POL" swrid="5626910" athleteid="5626910">
              <RESULTS>
                <RESULT eventid="3" points="440" swimtime="00:00:58.92" resultid="175810552" heatid="33" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="475" swimtime="00:00:27.87" resultid="175810551" heatid="117" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Makowski" birthdate="1987-01-13" gender="M" nation="POL" swrid="5626917" athleteid="5626917">
              <RESULTS>
                <RESULT eventid="3" points="295" swimtime="00:01:07.30" resultid="175810497" heatid="28" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="286" swimtime="00:00:37.84" resultid="175810495" heatid="87" lane="4" />
                <RESULT eventid="18" points="239" swimtime="00:01:29.04" resultid="175810498" heatid="96" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="226" swimtime="00:03:17.02" resultid="175810496" heatid="107" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                    <SPLIT distance="100" swimtime="00:01:30.08" />
                    <SPLIT distance="150" swimtime="00:02:22.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Krzekotowski" birthdate="1966-06-29" gender="M" nation="POL" swrid="5416779" athleteid="5416779">
              <RESULTS>
                <RESULT eventid="5" points="115" swimtime="00:03:23.91" resultid="175810245" heatid="44" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                    <SPLIT distance="100" swimtime="00:01:38.04" />
                    <SPLIT distance="150" swimtime="00:02:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="106" swimtime="00:07:28.08" resultid="175810248" heatid="54" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.19" />
                    <SPLIT distance="100" swimtime="00:01:44.18" />
                    <SPLIT distance="150" swimtime="00:02:40.63" />
                    <SPLIT distance="200" swimtime="00:04:36.10" />
                    <SPLIT distance="250" swimtime="00:06:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="58" swimtime="00:04:31.79" resultid="175810247" heatid="71" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.45" />
                    <SPLIT distance="100" swimtime="00:02:14.20" />
                    <SPLIT distance="150" swimtime="00:03:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" points="106" swimtime="00:03:51.50" resultid="175810246" heatid="133" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.45" />
                    <SPLIT distance="100" swimtime="00:01:59.00" />
                    <SPLIT distance="150" swimtime="00:02:59.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej Marek" lastname="Twarowski" birthdate="1965-05-24" gender="M" nation="POL" swrid="5125743" athleteid="5125743">
              <RESULTS>
                <RESULT eventid="5" points="147" swimtime="00:03:08.24" resultid="175810257" heatid="44" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                    <SPLIT distance="100" swimtime="00:01:33.77" />
                    <SPLIT distance="150" swimtime="00:02:23.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="157" swimtime="00:06:32.77" resultid="175810259" heatid="54" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.50" />
                    <SPLIT distance="100" swimtime="00:01:32.93" />
                    <SPLIT distance="150" swimtime="00:02:22.78" />
                    <SPLIT distance="200" swimtime="00:03:14.88" />
                    <SPLIT distance="250" swimtime="00:04:05.87" />
                    <SPLIT distance="300" swimtime="00:04:56.75" />
                    <SPLIT distance="350" swimtime="00:05:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11" points="163" swimtime="00:01:28.46" resultid="175810256" heatid="64" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="149" swimtime="00:03:19.18" resultid="175810258" heatid="71" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                    <SPLIT distance="100" swimtime="00:01:39.25" />
                    <SPLIT distance="150" swimtime="00:02:30.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Dusza" birthdate="1983-10-11" gender="F" nation="POL" swrid="5626902" athleteid="5626902">
              <RESULTS>
                <RESULT eventid="6" points="250" swimtime="00:02:54.94" resultid="175810314" heatid="45" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:23.23" />
                    <SPLIT distance="150" swimtime="00:02:09.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8" points="254" swimtime="00:06:08.92" resultid="175810315" heatid="53" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:12.16" />
                    <SPLIT distance="200" swimtime="00:03:00.00" />
                    <SPLIT distance="250" swimtime="00:03:47.69" />
                    <SPLIT distance="300" swimtime="00:04:35.36" />
                    <SPLIT distance="350" swimtime="00:05:23.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="27" points="219" swimtime="00:03:22.01" resultid="175810316" heatid="135" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                    <SPLIT distance="100" swimtime="00:01:39.28" />
                    <SPLIT distance="150" swimtime="00:02:36.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="208" swimtime="00:01:35.28" resultid="175810317" heatid="137" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Kubiak" birthdate="1989-07-05" gender="M" nation="POL" swrid="5626912" athleteid="5626912">
              <RESULTS>
                <RESULT eventid="5" points="232" swimtime="00:02:41.57" resultid="175810233" heatid="35" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="150" swimtime="00:02:00.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" points="120" swimtime="00:01:36.70" resultid="175810234" heatid="124" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Kular" birthdate="1987-08-28" gender="M" nation="POL" swrid="5626913" athleteid="5626913">
              <RESULTS>
                <RESULT eventid="5" points="189" swimtime="00:02:52.86" resultid="175810337" heatid="43" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                    <SPLIT distance="100" swimtime="00:01:20.46" />
                    <SPLIT distance="150" swimtime="00:02:06.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="180" swimtime="00:06:15.90" resultid="175810338" heatid="54" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:01:24.22" />
                    <SPLIT distance="150" swimtime="00:02:10.78" />
                    <SPLIT distance="200" swimtime="00:02:59.29" />
                    <SPLIT distance="250" swimtime="00:03:49.42" />
                    <SPLIT distance="300" swimtime="00:04:40.08" />
                    <SPLIT distance="350" swimtime="00:05:30.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Nechling" birthdate="1991-11-16" gender="F" nation="POL" swrid="5626923" athleteid="5626923">
              <RESULTS>
                <RESULT eventid="6" points="146" swimtime="00:03:29.40" resultid="175810255" heatid="38" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.57" />
                    <SPLIT distance="100" swimtime="00:01:37.70" />
                    <SPLIT distance="150" swimtime="00:02:33.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Grochowski" birthdate="1991-08-29" gender="M" nation="POL" swrid="5464090" athleteid="5464090">
              <RESULTS>
                <RESULT eventid="7" points="338" swimtime="00:05:04.50" resultid="175810282" heatid="48" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:50.64" />
                    <SPLIT distance="200" swimtime="00:02:29.13" />
                    <SPLIT distance="250" swimtime="00:03:07.53" />
                    <SPLIT distance="300" swimtime="00:03:46.34" />
                    <SPLIT distance="350" swimtime="00:04:24.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11" points="244" swimtime="00:01:17.29" resultid="175810279" heatid="66" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="254" swimtime="00:00:34.34" resultid="175810281" heatid="122" lane="3" />
                <RESULT eventid="24" points="213" swimtime="00:01:19.90" resultid="175810280" heatid="127" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kateryna" lastname="Moiseienko" birthdate="1979-12-22" gender="F" nation="POL" swrid="5484416" athleteid="5484416">
              <RESULTS>
                <RESULT eventid="8" points="82" swimtime="00:08:58.11" resultid="175810554" heatid="51" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.50" />
                    <SPLIT distance="100" swimtime="00:01:55.23" />
                    <SPLIT distance="150" swimtime="00:03:03.98" />
                    <SPLIT distance="200" swimtime="00:04:14.84" />
                    <SPLIT distance="250" swimtime="00:05:27.35" />
                    <SPLIT distance="300" swimtime="00:06:39.56" />
                    <SPLIT distance="350" swimtime="00:07:50.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="97" swimtime="00:04:18.18" resultid="175810553" heatid="76" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.81" />
                    <SPLIT distance="100" swimtime="00:02:02.92" />
                    <SPLIT distance="150" swimtime="00:03:11.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernard" lastname="Poloczek" birthdate="1947-02-25" gender="M" nation="POL" swrid="4792004" athleteid="4792004">
              <RESULTS>
                <RESULT eventid="9" points="122" swimtime="00:00:44.77" resultid="175810501" heatid="56" lane="3" />
                <RESULT eventid="11" points="111" swimtime="00:01:40.48" resultid="175810499" heatid="63" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="110" swimtime="00:00:45.36" resultid="175810500" heatid="115" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rudolf" lastname="Bugla" birthdate="1940-05-16" gender="M" nation="SVK" swrid="4831499" athleteid="4831499">
              <RESULTS>
                <RESULT eventid="9" points="18" swimtime="00:01:24.45" resultid="175810513" heatid="56" lane="4" />
                <RESULT eventid="16" points="30" swimtime="00:01:20.11" resultid="175810510" heatid="90" lane="5" />
                <RESULT eventid="18" points="34" swimtime="00:02:50.49" resultid="175810512" heatid="100" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="32" swimtime="00:06:16.05" resultid="175810511" heatid="104" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.56" />
                    <SPLIT distance="100" swimtime="00:03:04.30" />
                    <SPLIT distance="150" swimtime="00:04:40.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Ciecior" birthdate="1953-11-24" gender="M" nation="POL" swrid="4934027" athleteid="4934027">
              <RESULTS>
                <RESULT eventid="9" points="152" swimtime="00:00:41.56" resultid="175810509" heatid="57" lane="5" />
                <RESULT eventid="11" points="118" swimtime="00:01:38.29" resultid="175810506" heatid="63" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="123" swimtime="00:03:31.98" resultid="175810508" heatid="71" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.60" />
                    <SPLIT distance="100" swimtime="00:01:44.21" />
                    <SPLIT distance="150" swimtime="00:02:39.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" points="79" swimtime="00:01:50.92" resultid="175810507" heatid="124" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Dziedziczak-Szmytke" birthdate="1971-02-24" gender="F" nation="POL" swrid="5626903" athleteid="5626903">
              <RESULTS>
                <RESULT eventid="10" points="191" swimtime="00:00:43.84" resultid="175810285" heatid="62" lane="1" />
                <RESULT eventid="12" points="184" swimtime="00:01:36.34" resultid="175810283" heatid="68" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="189" swimtime="00:03:26.97" resultid="175810284" heatid="74" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                    <SPLIT distance="100" swimtime="00:01:38.01" />
                    <SPLIT distance="150" swimtime="00:02:32.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Wodyński" birthdate="1977-03-01" gender="M" nation="POL" swrid="5626946" athleteid="5626946">
              <RESULTS>
                <RESULT eventid="11" points="107" swimtime="00:01:41.75" resultid="175810562" heatid="64" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Radoslaw" lastname="Stefurak" birthdate="1974-09-07" gender="M" nation="POL" swrid="4429483" athleteid="4429483">
              <RESULTS>
                <RESULT eventid="16" points="283" swimtime="00:00:37.96" resultid="175810310" heatid="87" lane="2" />
                <RESULT eventid="18" points="272" swimtime="00:01:25.30" resultid="175810312" heatid="99" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="279" swimtime="00:03:03.71" resultid="175810311" heatid="110" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.87" />
                    <SPLIT distance="100" swimtime="00:01:26.23" />
                    <SPLIT distance="150" swimtime="00:02:13.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="218" swimtime="00:01:21.79" resultid="175810313" heatid="141" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Opałko" birthdate="1999-07-06" gender="F" nation="POL" swrid="4493246" athleteid="4493246">
              <RESULTS>
                <RESULT eventid="15" points="427" swimtime="00:00:37.91" resultid="175810514" heatid="80" lane="5" />
                <RESULT eventid="21" points="380" swimtime="00:00:33.65" resultid="175810516" heatid="118" lane="3" />
                <RESULT eventid="27" points="354" swimtime="00:02:52.14" resultid="175810515" heatid="131" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:18.13" />
                    <SPLIT distance="150" swimtime="00:02:08.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="398" swimtime="00:01:16.80" resultid="175810517" heatid="138" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Okaj" birthdate="2002-11-08" gender="F" nation="POL" swrid="4780566" athleteid="4780566">
              <RESULTS>
                <RESULT eventid="15" points="497" swimtime="00:00:36.04" resultid="175810327" heatid="88" lane="2" />
                <RESULT eventid="17" points="551" swimtime="00:01:16.04" resultid="175810329" heatid="101" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="27" points="480" swimtime="00:02:35.58" resultid="175810328" heatid="131" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:12.06" />
                    <SPLIT distance="150" swimtime="00:01:56.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="501" swimtime="00:01:11.12" resultid="175810330" heatid="146" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wieslaw" lastname="Majcher" birthdate="1950-09-19" gender="M" nation="POL" swrid="5240919" athleteid="5240919">
              <RESULTS>
                <RESULT eventid="16" points="40" swimtime="00:01:12.79" resultid="175810559" heatid="81" lane="2" />
                <RESULT eventid="18" points="36" swimtime="00:02:47.07" resultid="175810561" heatid="93" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="32" swimtime="00:06:18.28" resultid="175810560" heatid="104" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.81" />
                    <SPLIT distance="100" swimtime="00:02:57.03" />
                    <SPLIT distance="150" swimtime="00:04:37.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Krupiński" birthdate="1987-02-05" gender="M" nation="POL" swrid="5568771" athleteid="5568771">
              <RESULTS>
                <RESULT eventid="16" points="163" swimtime="00:00:45.67" resultid="175810529" heatid="79" lane="1" />
                <RESULT eventid="18" points="162" swimtime="00:01:41.33" resultid="175810531" heatid="94" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="163" swimtime="00:03:39.78" resultid="175810530" heatid="106" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                    <SPLIT distance="100" swimtime="00:01:42.52" />
                    <SPLIT distance="150" swimtime="00:02:40.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="166" swimtime="00:00:39.56" resultid="175810532" heatid="119" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Grzelczak" birthdate="1985-01-11" gender="M" nation="POL" swrid="5626906" athleteid="5626906">
              <RESULTS>
                <RESULT eventid="16" points="224" swimtime="00:00:41.04" resultid="175810275" heatid="82" lane="3" />
                <RESULT eventid="18" points="200" swimtime="00:01:34.42" resultid="175810278" heatid="94" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="180" swimtime="00:03:32.64" resultid="175810276" heatid="106" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.67" />
                    <SPLIT distance="100" swimtime="00:01:39.57" />
                    <SPLIT distance="150" swimtime="00:02:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="115" swimtime="00:00:44.62" resultid="175810277" heatid="115" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stefan" lastname="Niedzielski" birthdate="1955-02-13" gender="M" nation="POL" swrid="5626924" athleteid="5626924">
              <RESULTS>
                <RESULT eventid="16" points="115" swimtime="00:00:51.16" resultid="175810265" heatid="90" lane="2" />
                <RESULT eventid="18" points="113" swimtime="00:01:54.01" resultid="175810267" heatid="100" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="109" swimtime="00:04:11.34" resultid="175810266" heatid="106" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.64" />
                    <SPLIT distance="100" swimtime="00:01:59.49" />
                    <SPLIT distance="150" swimtime="00:03:05.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Szewczyk-Jachym" birthdate="1996-12-27" gender="M" nation="POL" swrid="5626938" athleteid="5626938">
              <RESULTS>
                <RESULT eventid="16" points="454" swimtime="00:00:32.45" resultid="175810271" heatid="89" lane="6" />
                <RESULT eventid="18" points="423" swimtime="00:01:13.63" resultid="175810274" heatid="95" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="421" swimtime="00:00:29.00" resultid="175810273" heatid="117" lane="6" />
                <RESULT eventid="24" points="360" swimtime="00:01:07.13" resultid="175810272" heatid="126" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Galon" birthdate="1995-05-21" gender="M" nation="POL" swrid="4265580" athleteid="4265580">
              <RESULTS>
                <RESULT eventid="28" points="555" swimtime="00:02:13.39" resultid="175810260" heatid="136" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.86" />
                    <SPLIT distance="100" swimtime="00:01:01.33" />
                    <SPLIT distance="150" swimtime="00:01:39.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="31" points="255" swimtime="00:02:18.58" resultid="175810304" heatid="149" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="150" swimtime="00:01:49.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5468089" number="1" />
                    <RELAYPOSITION athleteid="5626926" number="2" />
                    <RELAYPOSITION athleteid="5484408" number="3" />
                    <RELAYPOSITION athleteid="5626897" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="31" points="257" swimtime="00:02:18.07" resultid="175810325" heatid="149" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:07.47" />
                    <SPLIT distance="150" swimtime="00:01:44.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5626895" number="1" />
                    <RELAYPOSITION athleteid="5626920" number="2" />
                    <RELAYPOSITION athleteid="5626902" number="3" />
                    <RELAYPOSITION athleteid="4429483" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="198" swimtime="00:02:44.93" resultid="175810305" heatid="153" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5626926" number="1" />
                    <RELAYPOSITION athleteid="5468089" number="2" />
                    <RELAYPOSITION athleteid="5626897" number="3" />
                    <RELAYPOSITION athleteid="5484408" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="218" swimtime="00:02:39.70" resultid="175810326" heatid="153" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.05" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="150" swimtime="00:02:06.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5626895" number="1" />
                    <RELAYPOSITION athleteid="4429483" number="2" />
                    <RELAYPOSITION athleteid="5626902" number="3" />
                    <RELAYPOSITION athleteid="5626920" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02211" nation="POL" region="11" clubid="85535" swrid="85535" name="MUKS Gilus Gilowice">
          <ATHLETES>
            <ATHLETE firstname="Sławomir" lastname="Formas" birthdate="1969-11-05" gender="M" nation="POL" license="502211700187" swrid="4292540" athleteid="4292540">
              <RESULTS>
                <RESULT eventid="16" points="514" swimtime="00:00:31.13" resultid="175810585" heatid="89" lane="4" />
                <RESULT eventid="18" points="519" swimtime="00:01:08.77" resultid="175810587" heatid="95" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="494" swimtime="00:02:31.95" resultid="175810586" heatid="105" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                    <SPLIT distance="150" swimtime="00:01:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="425" swimtime="00:01:05.54" resultid="175810588" heatid="142" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03415" nation="POL" region="15" clubid="86514" swrid="86514" name="Uczniowski Klub Sportowy City Zen Poznań" shortname="UKS City Zen Poznań">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Lutowicz" birthdate="1950-08-23" gender="F" nation="POL" swrid="4188428" athleteid="4188428">
              <RESULTS>
                <RESULT eventid="2" points="84" swimtime="00:00:52.34" resultid="175810389" heatid="16" lane="4" />
                <RESULT eventid="10" points="80" swimtime="00:00:58.58" resultid="175810390" heatid="61" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Matyszczak" birthdate="1970-12-14" gender="M" nation="POL" swrid="5471729" athleteid="5471729">
              <RESULTS>
                <RESULT eventid="1" points="282" swimtime="00:00:30.71" resultid="175810395" heatid="6" lane="3" />
                <RESULT eventid="3" points="254" swimtime="00:01:10.73" resultid="175810397" heatid="24" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="225" swimtime="00:02:43.19" resultid="175810396" heatid="35" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:17.70" />
                    <SPLIT distance="150" swimtime="00:02:00.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="182" swimtime="00:01:26.92" resultid="175810398" heatid="144" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Pietraszewski" birthdate="1955-04-07" gender="M" nation="POL" swrid="4187282" athleteid="4187282">
              <RESULTS>
                <RESULT eventid="1" points="104" swimtime="00:00:42.83" resultid="175810399" heatid="14" lane="1" />
                <RESULT eventid="3" points="114" swimtime="00:01:32.33" resultid="175810401" heatid="31" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="68" swimtime="00:00:54.21" resultid="175810402" heatid="56" lane="6" />
                <RESULT eventid="11" points="66" swimtime="00:01:59.52" resultid="175810400" heatid="63" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Rolewski" birthdate="1967-01-01" gender="M" nation="POL" swrid="5626933" athleteid="5626933">
              <RESULTS>
                <RESULT eventid="1" points="17" swimtime="00:01:17.97" resultid="175810417" heatid="3" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rusłana" lastname="Dembecka" birthdate="1957-10-01" gender="F" nation="POL" swrid="5626901" athleteid="5626901">
              <RESULTS>
                <RESULT eventid="10" points="56" swimtime="00:01:05.76" resultid="175810416" heatid="61" lane="2" />
                <RESULT eventid="15" points="119" swimtime="00:00:57.99" resultid="175810413" heatid="86" lane="2" />
                <RESULT eventid="17" points="107" swimtime="00:02:10.98" resultid="175810415" heatid="97" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="111" swimtime="00:04:39.86" resultid="175810414" heatid="108" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.03" />
                    <SPLIT distance="100" swimtime="00:02:15.53" />
                    <SPLIT distance="150" swimtime="00:03:28.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Łasińska-Błachowicz" birthdate="1954-07-13" gender="F" nation="POL" swrid="5471727" athleteid="5471727">
              <RESULTS>
                <RESULT eventid="12" points="68" swimtime="00:02:14.43" resultid="175810405" heatid="69" lane="5" />
                <RESULT eventid="21" points="57" swimtime="00:01:03.00" resultid="175810407" heatid="118" lane="6" />
                <RESULT eventid="27" points="72" swimtime="00:04:52.15" resultid="175810406" heatid="135" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.30" />
                    <SPLIT distance="100" swimtime="00:02:25.93" />
                    <SPLIT distance="150" swimtime="00:03:42.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="82" swimtime="00:02:09.98" resultid="175810408" heatid="143" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Slawomir" lastname="Cybertowicz" birthdate="1966-01-12" gender="M" nation="POL" swrid="4269915" athleteid="4269915">
              <RESULTS>
                <RESULT eventid="16" points="240" swimtime="00:00:40.11" resultid="175810403" heatid="83" lane="5" />
                <RESULT eventid="18" points="233" swimtime="00:01:29.82" resultid="175810404" heatid="99" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Rybak-Starczak" birthdate="1975-01-16" gender="F" nation="POL" swrid="5439532" athleteid="5439532">
              <RESULTS>
                <RESULT eventid="17" points="309" swimtime="00:01:32.22" resultid="175810393" heatid="98" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="308" swimtime="00:03:19.24" resultid="175810392" heatid="112" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                    <SPLIT distance="100" swimtime="00:01:36.91" />
                    <SPLIT distance="150" swimtime="00:02:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="27" points="271" status="DSQ" swimtime="00:03:08.22" resultid="175810391" heatid="131" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:01:33.17" />
                    <SPLIT distance="150" swimtime="00:02:24.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="281" swimtime="00:01:26.19" resultid="175810394" heatid="137" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Putowska" birthdate="1962-01-22" gender="F" nation="POL" swrid="5416834" athleteid="5416834">
              <RESULTS>
                <RESULT eventid="17" points="174" swimtime="00:01:51.66" resultid="175810411" heatid="98" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="183" swimtime="00:03:57.02" resultid="175810410" heatid="109" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.30" />
                    <SPLIT distance="100" swimtime="00:01:52.98" />
                    <SPLIT distance="150" swimtime="00:02:56.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="26" points="82" swimtime="00:04:34.90" resultid="175810412" heatid="129" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.37" />
                    <SPLIT distance="100" swimtime="00:02:04.73" />
                    <SPLIT distance="150" swimtime="00:03:21.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="27" points="124" swimtime="00:04:03.74" resultid="175810409" heatid="135" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.94" />
                    <SPLIT distance="100" swimtime="00:02:00.24" />
                    <SPLIT distance="150" swimtime="00:03:04.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="31" points="126" swimtime="00:02:55.08" resultid="175810418" heatid="148" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.44" />
                    <SPLIT distance="100" swimtime="00:01:31.29" />
                    <SPLIT distance="150" swimtime="00:02:24.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5471727" number="1" />
                    <RELAYPOSITION athleteid="4187282" number="2" />
                    <RELAYPOSITION athleteid="5626901" number="3" />
                    <RELAYPOSITION athleteid="5471729" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="183" swimtime="00:02:49.36" resultid="175810419" heatid="151" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                    <SPLIT distance="100" swimtime="00:01:23.22" />
                    <SPLIT distance="150" swimtime="00:02:15.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5471729" number="1" />
                    <RELAYPOSITION athleteid="5439532" number="2" />
                    <RELAYPOSITION athleteid="5416834" number="3" />
                    <RELAYPOSITION athleteid="4269915" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03508" nation="POL" region="08" clubid="79441" swrid="79441" name="KS PRESTIGE Rzeszów">
          <ATHLETES>
            <ATHLETE firstname="Patrycja" lastname="Rupa" birthdate="1996-01-11" gender="F" nation="POL" license="103508600006" swrid="4108567" athleteid="4108567">
              <RESULTS>
                <RESULT eventid="10" points="453" swimtime="00:00:32.88" resultid="175810423" heatid="62" lane="2" />
                <RESULT eventid="12" points="456" swimtime="00:01:11.28" resultid="175810420" heatid="68" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="416" swimtime="00:02:39.28" resultid="175810422" heatid="76" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:17.70" />
                    <SPLIT distance="150" swimtime="00:01:58.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="280" swimtime="00:03:25.51" resultid="175810421" heatid="102" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.08" />
                    <SPLIT distance="100" swimtime="00:01:40.15" />
                    <SPLIT distance="150" swimtime="00:02:32.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02805" nation="POL" region="05" clubid="86339" swrid="86339" name="MUKS Zgierz">
          <ATHLETES>
            <ATHLETE firstname="Urszula" lastname="Mróz" birthdate="1962-03-03" gender="F" nation="POL" license="502805600024" swrid="4754660" athleteid="4754660">
              <RESULTS>
                <RESULT eventid="2" points="313" swimtime="00:00:33.75" resultid="175809862" heatid="4" lane="6" />
                <RESULT eventid="4" points="291" swimtime="00:01:15.78" resultid="175809864" heatid="22" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" points="261" swimtime="00:00:44.66" resultid="175809863" heatid="80" lane="6" />
                <RESULT eventid="29" points="295" swimtime="00:01:24.83" resultid="175809865" heatid="137" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Rembowska-Świeboda" birthdate="1968-06-27" gender="F" nation="POL" swrid="5439505" athleteid="5439505">
              <RESULTS>
                <RESULT eventid="2" points="318" swimtime="00:00:33.57" resultid="175809873" heatid="5" lane="3" />
                <RESULT eventid="4" points="285" swimtime="00:01:16.32" resultid="175809875" heatid="23" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10" points="296" swimtime="00:00:37.88" resultid="175809876" heatid="58" lane="5" />
                <RESULT eventid="12" points="284" swimtime="00:01:23.43" resultid="175809874" heatid="65" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Przytulski" birthdate="1957-01-09" gender="M" nation="POL" license="502805700049" swrid="4754657" athleteid="4754657">
              <RESULTS>
                <RESULT eventid="1" points="240" swimtime="00:00:32.40" resultid="175809896" heatid="6" lane="1" />
                <RESULT eventid="22" points="253" swimtime="00:00:34.37" resultid="175809898" heatid="114" lane="2" />
                <RESULT eventid="28" points="210" swimtime="00:03:04.34" resultid="175809897" heatid="132" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:26.56" />
                    <SPLIT distance="150" swimtime="00:02:24.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="217" swimtime="00:01:21.94" resultid="175809899" heatid="140" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisław" lastname="Jasiński" birthdate="1960-07-23" gender="M" nation="POL" license="502805700027" swrid="5374015" athleteid="5374015">
              <RESULTS>
                <RESULT eventid="1" points="209" swimtime="00:00:33.93" resultid="175809900" heatid="7" lane="5" />
                <RESULT eventid="3" points="187" swimtime="00:01:18.29" resultid="175809902" heatid="25" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" points="132" swimtime="00:03:35.29" resultid="175809901" heatid="133" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.43" />
                    <SPLIT distance="100" swimtime="00:01:47.68" />
                    <SPLIT distance="150" swimtime="00:02:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="139" status="DSQ" swimtime="00:01:35.03" resultid="175809903" heatid="141" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Gołębiowski" birthdate="1996-09-02" gender="M" nation="POL" swrid="4115580" athleteid="4115580">
              <RESULTS>
                <RESULT eventid="1" points="425" swimtime="00:00:26.81" resultid="175809904" heatid="8" lane="6" />
                <RESULT eventid="9" points="373" swimtime="00:00:30.85" resultid="175809907" heatid="59" lane="1" />
                <RESULT eventid="16" points="388" swimtime="00:00:34.18" resultid="175809905" heatid="84" lane="5" />
                <RESULT eventid="18" points="416" swimtime="00:01:14.03" resultid="175809906" heatid="96" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Węgrzycka" birthdate="1977-01-26" gender="F" nation="POL" license="502805600056" swrid="5464095" athleteid="5464095">
              <RESULTS>
                <RESULT eventid="2" points="177" swimtime="00:00:40.79" resultid="175809912" heatid="9" lane="1" />
                <RESULT eventid="4" points="147" swimtime="00:01:35.16" resultid="175809914" heatid="26" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" points="147" status="DSQ" swimtime="00:00:54.07" resultid="175809913" heatid="85" lane="1" />
                <RESULT eventid="17" points="132" swimtime="00:02:02.33" resultid="175809915" heatid="97" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Ścibiorek" birthdate="1997-02-19" gender="M" nation="POL" swrid="4287843" athleteid="4287843">
              <RESULTS>
                <RESULT eventid="1" points="462" swimtime="00:00:26.07" resultid="175809920" heatid="8" lane="1" />
                <RESULT eventid="11" points="372" swimtime="00:01:07.14" resultid="175809921" heatid="66" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="440" swimtime="00:00:28.58" resultid="175809922" heatid="117" lane="1" />
                <RESULT eventid="30" points="416" swimtime="00:01:06.01" resultid="175809923" heatid="142" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Ławniczak" birthdate="1979-09-13" gender="F" nation="POL" swrid="5626914" athleteid="5626914">
              <RESULTS>
                <RESULT eventid="2" points="201" swimtime="00:00:39.10" resultid="175809928" heatid="10" lane="4" />
                <RESULT eventid="4" points="165" swimtime="00:01:31.46" resultid="175809930" heatid="27" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" points="209" swimtime="00:00:48.08" resultid="175809929" heatid="78" lane="5" />
                <RESULT eventid="29" points="161" swimtime="00:01:43.70" resultid="175809931" heatid="143" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Pietruszewski - Gil" birthdate="1986-12-17" gender="M" nation="POL" swrid="5626930" athleteid="5626930">
              <RESULTS>
                <RESULT eventid="1" points="266" swimtime="00:00:31.33" resultid="175809932" heatid="2" lane="2" />
                <RESULT eventid="3" points="263" swimtime="00:01:09.97" resultid="175809934" heatid="28" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="187" swimtime="00:00:43.57" resultid="175809933" heatid="82" lane="1" />
                <RESULT eventid="30" points="208" swimtime="00:01:23.16" resultid="175809935" heatid="144" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dagmara" lastname="Luzniakowska" birthdate="1980-04-29" gender="F" nation="POL" swrid="5582458" athleteid="5582458">
              <RESULTS>
                <RESULT eventid="2" points="225" swimtime="00:00:37.65" resultid="175809940" heatid="10" lane="5" />
                <RESULT eventid="4" points="212" swimtime="00:01:24.22" resultid="175809943" heatid="22" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" points="258" swimtime="00:02:53.16" resultid="175809941" heatid="38" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:23.62" />
                    <SPLIT distance="150" swimtime="00:02:09.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" points="183" swimtime="00:00:42.87" resultid="175809942" heatid="118" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Morozowski" birthdate="1973-05-09" gender="M" nation="POL" license="102805700051" swrid="5416829" athleteid="5416829">
              <RESULTS>
                <RESULT eventid="3" points="238" swimtime="00:01:12.34" resultid="175809886" heatid="24" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="195" swimtime="00:06:05.49" resultid="175809887" heatid="47" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="150" swimtime="00:02:05.81" />
                    <SPLIT distance="200" swimtime="00:02:52.70" />
                    <SPLIT distance="250" swimtime="00:03:41.22" />
                    <SPLIT distance="300" swimtime="00:04:30.68" />
                    <SPLIT distance="350" swimtime="00:05:19.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="255" swimtime="00:00:39.30" resultid="175809884" heatid="83" lane="3" />
                <RESULT eventid="20" points="185" swimtime="00:03:30.56" resultid="175809885" heatid="106" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.33" />
                    <SPLIT distance="100" swimtime="00:01:40.44" />
                    <SPLIT distance="150" swimtime="00:02:35.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Dziedziczak" birthdate="1977-02-04" gender="M" nation="POL" swrid="5558378" athleteid="5558378">
              <RESULTS>
                <RESULT eventid="3" points="261" swimtime="00:01:10.15" resultid="175809894" heatid="24" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="189" swimtime="00:06:09.76" resultid="175809895" heatid="48" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:20.03" />
                    <SPLIT distance="150" swimtime="00:02:05.90" />
                    <SPLIT distance="200" swimtime="00:02:54.48" />
                    <SPLIT distance="250" swimtime="00:03:43.84" />
                    <SPLIT distance="300" swimtime="00:04:34.70" />
                    <SPLIT distance="350" swimtime="00:05:24.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11" points="168" swimtime="00:01:27.46" resultid="175809892" heatid="66" lane="3" />
                <RESULT eventid="28" points="212" swimtime="00:03:03.62" resultid="175809893" heatid="132" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:25.60" />
                    <SPLIT distance="150" swimtime="00:02:24.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="503605600029" swrid="5464091" athleteid="5464091">
              <RESULTS>
                <RESULT eventid="8" points="180" swimtime="00:06:54.27" resultid="175809947" heatid="49" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                    <SPLIT distance="100" swimtime="00:01:34.60" />
                    <SPLIT distance="150" swimtime="00:02:27.77" />
                    <SPLIT distance="200" swimtime="00:03:21.20" />
                    <SPLIT distance="250" swimtime="00:04:15.05" />
                    <SPLIT distance="300" swimtime="00:05:08.64" />
                    <SPLIT distance="350" swimtime="00:06:03.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="185" swimtime="00:03:56.14" resultid="175809945" heatid="109" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.09" />
                    <SPLIT distance="100" swimtime="00:01:54.77" />
                    <SPLIT distance="150" swimtime="00:02:55.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="26" points="124" swimtime="00:03:59.33" resultid="175809946" heatid="129" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.80" />
                    <SPLIT distance="100" swimtime="00:01:53.28" />
                    <SPLIT distance="150" swimtime="00:02:56.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="27" points="157" swimtime="00:03:45.48" resultid="175809944" heatid="135" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.26" />
                    <SPLIT distance="100" swimtime="00:01:51.67" />
                    <SPLIT distance="150" swimtime="00:02:55.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Sypniewski" birthdate="1957-01-02" gender="M" nation="POL" swrid="5373999" athleteid="5373999">
              <RESULTS>
                <RESULT eventid="9" points="175" swimtime="00:00:39.67" resultid="175809869" heatid="57" lane="4" />
                <RESULT eventid="11" points="163" swimtime="00:01:28.47" resultid="175809866" heatid="64" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="191" swimtime="00:00:43.30" resultid="175809867" heatid="81" lane="3" />
                <RESULT eventid="18" points="187" swimtime="00:01:36.54" resultid="175809868" heatid="94" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Matczak" birthdate="1989-08-12" gender="M" nation="POL" swrid="4071609" athleteid="4071609">
              <RESULTS>
                <RESULT eventid="11" points="439" swimtime="00:01:03.55" resultid="175809881" heatid="66" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" points="523" swimtime="00:01:08.57" resultid="175809883" heatid="95" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="556" swimtime="00:02:26.07" resultid="175809882" heatid="105" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="150" swimtime="00:01:47.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Wiczel" birthdate="1948-01-22" gender="M" nation="POL" swrid="4876444" athleteid="4876444">
              <RESULTS>
                <RESULT eventid="13" points="108" swimtime="00:03:41.40" resultid="175809891" heatid="71" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.22" />
                    <SPLIT distance="100" swimtime="00:01:50.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="180" swimtime="00:00:44.15" resultid="175809888" heatid="82" lane="6" />
                <RESULT eventid="18" points="178" swimtime="00:01:38.25" resultid="175809890" heatid="94" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="167" swimtime="00:03:38.05" resultid="175809889" heatid="106" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.56" />
                    <SPLIT distance="100" swimtime="00:01:46.57" />
                    <SPLIT distance="150" swimtime="00:02:44.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Wypych - Staszewska" birthdate="1970-08-16" gender="F" nation="POL" swrid="5626948" athleteid="5626948">
              <RESULTS>
                <RESULT eventid="14" points="187" swimtime="00:03:27.68" resultid="175809938" heatid="72" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.18" />
                    <SPLIT distance="100" swimtime="00:01:41.83" />
                    <SPLIT distance="150" swimtime="00:02:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" points="205" swimtime="00:01:32.46" resultid="175809937" heatid="123" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="26" points="182" swimtime="00:03:30.90" resultid="175809939" heatid="129" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:40.34" />
                    <SPLIT distance="150" swimtime="00:02:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="27" points="213" swimtime="00:03:23.75" resultid="175809936" heatid="134" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:01:36.63" />
                    <SPLIT distance="150" swimtime="00:02:38.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Woźniak" birthdate="1980-09-30" gender="M" nation="POL" swrid="5506643" athleteid="5506643">
              <RESULTS>
                <RESULT eventid="16" points="240" swimtime="00:00:40.10" resultid="175809877" heatid="82" lane="4" />
                <RESULT eventid="18" points="221" swimtime="00:01:31.32" resultid="175809879" heatid="94" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="207" swimtime="00:03:23.12" resultid="175809878" heatid="104" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:34.69" />
                    <SPLIT distance="150" swimtime="00:02:29.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="175" swimtime="00:01:27.98" resultid="175809880" heatid="139" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michal" lastname="Rudzinski" birthdate="1966-05-10" gender="M" nation="POL" license="510414700010" swrid="4934041" athleteid="4934041">
              <RESULTS>
                <RESULT eventid="16" points="168" swimtime="00:00:45.16" resultid="175809908" heatid="82" lane="5" />
                <RESULT eventid="20" points="171" swimtime="00:03:36.26" resultid="175809909" heatid="107" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.11" />
                    <SPLIT distance="100" swimtime="00:01:42.06" />
                    <SPLIT distance="150" swimtime="00:02:40.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="120" swimtime="00:00:44.09" resultid="175809910" heatid="115" lane="3" />
                <RESULT eventid="25" points="91" swimtime="00:04:00.05" resultid="175809911" heatid="128" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.18" />
                    <SPLIT distance="100" swimtime="00:01:49.64" />
                    <SPLIT distance="150" swimtime="00:02:54.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Wiśniewska" birthdate="1981-02-26" gender="F" nation="POL" license="502805600123" swrid="5464096" athleteid="5464096">
              <RESULTS>
                <RESULT eventid="15" points="131" swimtime="00:00:56.19" resultid="175809916" heatid="86" lane="1" />
                <RESULT eventid="17" points="116" swimtime="00:02:07.65" resultid="175809919" heatid="97" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="121" swimtime="00:04:31.80" resultid="175809917" heatid="108" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.69" />
                    <SPLIT distance="100" swimtime="00:02:10.13" />
                    <SPLIT distance="150" swimtime="00:03:22.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" points="79" swimtime="00:00:56.76" resultid="175809918" heatid="116" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1977-01-05" gender="F" nation="POL" license="502805600055" swrid="4655158" athleteid="4655158">
              <RESULTS>
                <RESULT eventid="15" points="234" swimtime="00:00:46.32" resultid="175809924" heatid="85" lane="3" />
                <RESULT eventid="17" points="229" swimtime="00:01:41.83" resultid="175809926" heatid="98" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="232" swimtime="00:03:38.91" resultid="175809925" heatid="109" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.01" />
                    <SPLIT distance="100" swimtime="00:01:46.76" />
                    <SPLIT distance="150" swimtime="00:02:42.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="170" swimtime="00:01:41.85" resultid="175809927" heatid="137" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Ścibiorek" birthdate="1971-09-12" gender="F" nation="POL" license="502805600026" swrid="4992745" athleteid="4992745">
              <RESULTS>
                <RESULT eventid="21" points="405" swimtime="00:00:32.94" resultid="175809871" heatid="113" lane="5" />
                <RESULT eventid="27" points="408" swimtime="00:02:44.21" resultid="175809870" heatid="131" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:16.38" />
                    <SPLIT distance="150" swimtime="00:02:04.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="412" swimtime="00:01:15.90" resultid="175809872" heatid="138" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="31" points="312" swimtime="00:02:09.47" resultid="175809948" heatid="149" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:04.26" />
                    <SPLIT distance="150" swimtime="00:01:37.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4992745" number="1" />
                    <RELAYPOSITION athleteid="5374015" number="2" />
                    <RELAYPOSITION athleteid="4754660" number="3" />
                    <RELAYPOSITION athleteid="4754657" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="31" points="271" swimtime="00:02:15.73" resultid="175809950" heatid="148" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:05.24" />
                    <SPLIT distance="150" swimtime="00:01:42.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5373999" number="1" />
                    <RELAYPOSITION athleteid="5439505" number="2" />
                    <RELAYPOSITION athleteid="5582458" number="3" />
                    <RELAYPOSITION athleteid="5416829" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="31" points="276" swimtime="00:02:14.98" resultid="175809952" heatid="149" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                    <SPLIT distance="150" swimtime="00:01:49.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5558378" number="1" />
                    <RELAYPOSITION athleteid="4655158" number="2" />
                    <RELAYPOSITION athleteid="5626914" number="3" />
                    <RELAYPOSITION athleteid="4287843" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="251" swimtime="00:02:32.44" resultid="175809949" heatid="151" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:01:20.74" />
                    <SPLIT distance="150" swimtime="00:02:00.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5439505" number="1" />
                    <RELAYPOSITION athleteid="5373999" number="2" />
                    <RELAYPOSITION athleteid="5626948" number="3" />
                    <RELAYPOSITION athleteid="4754657" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="216" swimtime="00:02:40.14" resultid="175809951" heatid="153" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:17.89" />
                    <SPLIT distance="150" swimtime="00:02:01.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4992745" number="1" />
                    <RELAYPOSITION athleteid="5416829" number="2" />
                    <RELAYPOSITION athleteid="4934041" number="3" />
                    <RELAYPOSITION athleteid="5582458" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="245" swimtime="00:02:33.52" resultid="175809953" heatid="153" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                    <SPLIT distance="100" swimtime="00:01:24.74" />
                    <SPLIT distance="150" swimtime="00:01:54.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5558378" number="1" />
                    <RELAYPOSITION athleteid="4655158" number="2" />
                    <RELAYPOSITION athleteid="4287843" number="3" />
                    <RELAYPOSITION athleteid="5626914" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="05215" nation="POL" region="15" clubid="90691" swrid="90691" name="MUKS HURAGAN Koło">
          <ATHLETES>
            <ATHLETE firstname="Joanna" lastname="Wojnicka" birthdate="1994-01-06" gender="F" nation="POL" swrid="5626947" athleteid="5626947">
              <RESULTS>
                <RESULT eventid="2" points="268" swimtime="00:00:35.55" resultid="175809958" heatid="10" lane="2" />
                <RESULT eventid="4" points="255" swimtime="00:01:19.18" resultid="175809960" heatid="27" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" points="234" swimtime="00:00:46.29" resultid="175809959" heatid="77" lane="3" />
                <RESULT eventid="17" points="211" swimtime="00:01:44.63" resultid="175809961" heatid="92" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PKMTR" nation="SVK" region="SSO" clubid="89401" swrid="89401" name="Plavecký klub Masters Turčianski raci" shortname="PKM Turčianski raci">
          <ATHLETES>
            <ATHLETE firstname="Katarína" lastname="Turanská" birthdate="1972-06-16" gender="F" nation="SVK" license="SVK17844" swrid="5101530" athleteid="5101530">
              <RESULTS>
                <RESULT eventid="2" points="108" swimtime="00:00:48.11" resultid="175810081" heatid="16" lane="3" />
                <RESULT eventid="15" points="193" swimtime="00:00:49.40" resultid="175810082" heatid="85" lane="5" />
                <RESULT eventid="19" points="163" swimtime="00:04:06.22" resultid="175810083" heatid="109" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.72" />
                    <SPLIT distance="100" swimtime="00:01:59.16" />
                    <SPLIT distance="150" swimtime="00:03:02.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Branislav" lastname="Turanský" birthdate="1967-12-18" gender="M" nation="SVK" license="SVK13190" swrid="4826051" athleteid="4826051">
              <RESULTS>
                <RESULT eventid="1" points="352" swimtime="00:00:28.55" resultid="175810084" heatid="18" lane="5" />
                <RESULT eventid="24" points="256" swimtime="00:01:15.16" resultid="175810085" heatid="126" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ján" lastname="Vanko" birthdate="1955-06-08" gender="M" nation="SVK" license="SVK17842" swrid="5101534" athleteid="5101534">
              <RESULTS>
                <RESULT eventid="1" points="190" swimtime="00:00:35.05" resultid="175810086" heatid="11" lane="2" />
                <RESULT eventid="16" points="147" swimtime="00:00:47.18" resultid="175810087" heatid="79" lane="3" />
                <RESULT eventid="28" points="124" swimtime="00:03:39.34" resultid="175810088" heatid="133" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.70" />
                    <SPLIT distance="100" swimtime="00:01:44.97" />
                    <SPLIT distance="150" swimtime="00:02:51.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04901" nation="POL" region="01" clubid="89936" swrid="89936" name="Klub Sportowy Neptun Świdnica" shortname="KS Neptun Świdnica">
          <ATHLETES>
            <ATHLETE firstname="Bartłomiej" lastname="Żukowski" birthdate="1993-04-26" gender="M" nation="POL" license="104901700097" swrid="4087259" athleteid="4087259">
              <RESULTS>
                <RESULT eventid="16" points="638" swimtime="00:00:28.97" resultid="175810424" heatid="89" lane="3" />
                <RESULT eventid="18" points="644" swimtime="00:01:03.99" resultid="175810426" heatid="95" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="585" swimtime="00:02:23.63" resultid="175810425" heatid="103" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="150" swimtime="00:01:46.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00612" nation="POL" region="12" clubid="65776" swrid="65776" name="KS KSZO Ostrowiec Świetokrzyski" shortname="KSZO Ostrowiec Świętokrzyski">
          <ATHLETES>
            <ATHLETE firstname="Stanisław" lastname="Sejmicki" birthdate="1961-05-04" gender="M" nation="POL" swrid="5558380" athleteid="5558380">
              <RESULTS>
                <RESULT eventid="1" points="162" swimtime="00:00:36.93" resultid="175810137" heatid="11" lane="6" />
                <RESULT eventid="16" points="197" swimtime="00:00:42.85" resultid="175810138" heatid="79" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="65887" swrid="65887" name="UKP UNIA Oświęcim">
          <ATHLETES>
            <ATHLETE firstname="Ilona" lastname="Szkudlarz" birthdate="1966-05-03" gender="F" nation="POL" swrid="4992932" athleteid="4992932">
              <RESULTS>
                <RESULT eventid="2" points="265" swimtime="00:00:35.68" resultid="175810223" heatid="10" lane="3" />
                <RESULT eventid="4" points="212" swimtime="00:01:24.20" resultid="175810225" heatid="27" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10" points="187" swimtime="00:00:44.16" resultid="175810227" heatid="62" lane="5" />
                <RESULT eventid="15" points="214" swimtime="00:00:47.73" resultid="175810224" heatid="78" lane="4" />
                <RESULT eventid="17" points="212" swimtime="00:01:44.57" resultid="175810226" heatid="92" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Lipniarska-Skubis" birthdate="1952-07-01" gender="F" nation="POL" swrid="5582457" athleteid="5582457">
              <RESULTS>
                <RESULT eventid="6" points="63" swimtime="00:04:36.08" resultid="175810231" heatid="38" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.20" />
                    <SPLIT distance="100" swimtime="00:02:12.53" />
                    <SPLIT distance="150" swimtime="00:03:24.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="76" swimtime="00:05:17.04" resultid="175810232" heatid="111" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.80" />
                    <SPLIT distance="100" swimtime="00:02:34.46" />
                    <SPLIT distance="150" swimtime="00:03:56.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jolanta" lastname="Płatek" birthdate="1971-09-10" gender="F" nation="POL" swrid="4992931" athleteid="4992931">
              <RESULTS>
                <RESULT eventid="10" points="262" swimtime="00:00:39.49" resultid="175810222" heatid="62" lane="4" />
                <RESULT eventid="12" points="239" swimtime="00:01:28.39" resultid="175810220" heatid="68" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="240" swimtime="00:03:11.37" resultid="175810221" heatid="76" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                    <SPLIT distance="100" swimtime="00:01:32.72" />
                    <SPLIT distance="150" swimtime="00:02:22.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Dorywalski" birthdate="1961-03-16" gender="M" nation="POL" swrid="4992929" athleteid="4992929">
              <RESULTS>
                <RESULT eventid="9" points="179" swimtime="00:00:39.42" resultid="175810230" heatid="60" lane="3" />
                <RESULT eventid="11" points="186" swimtime="00:01:24.55" resultid="175810228" heatid="66" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="187" swimtime="00:03:04.71" resultid="175810229" heatid="75" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                    <SPLIT distance="100" swimtime="00:01:29.17" />
                    <SPLIT distance="150" swimtime="00:02:17.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="NATION" code="UKR" nation="UKR" clubid="375" swrid="375" name="Ukraine">
          <ATHLETES>
            <ATHLETE firstname="Sergei" firstname.en="Serhii" lastname="Chernov" birthdate="1950-07-15" gender="M" nation="UKR" swrid="5610693" athleteid="5610693">
              <RESULTS>
                <RESULT eventid="1" points="46" swimtime="00:00:55.97" resultid="175810607" heatid="3" lane="3" />
                <RESULT eventid="3" points="37" swimtime="00:02:14.06" resultid="175810609" heatid="31" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="47" swimtime="00:04:34.76" resultid="175810608" heatid="40" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.82" />
                    <SPLIT distance="100" swimtime="00:02:12.31" />
                    <SPLIT distance="150" swimtime="00:03:24.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12914" nation="POL" region="14" clubid="83593" swrid="83593" name="Water Squad">
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Kaczmarek" birthdate="1985-05-07" gender="F" nation="POL" swrid="5240932" athleteid="5240932">
              <RESULTS>
                <RESULT eventid="2" points="419" swimtime="00:00:30.64" resultid="175810149" heatid="15" lane="6" />
                <RESULT eventid="10" points="458" swimtime="00:00:32.76" resultid="175810152" heatid="58" lane="3" />
                <RESULT eventid="27" points="433" swimtime="00:02:41.07" resultid="175810150" heatid="131" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:13.67" />
                    <SPLIT distance="150" swimtime="00:02:00.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="456" swimtime="00:01:13.41" resultid="175810151" heatid="138" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aneta" lastname="Dolińska" birthdate="1990-03-12" gender="F" nation="POL" swrid="4251116" athleteid="4251116">
              <RESULTS>
                <RESULT eventid="2" points="368" swimtime="00:00:31.97" resultid="175810153" heatid="4" lane="5" />
                <RESULT eventid="8" points="290" swimtime="00:05:53.37" resultid="175810156" heatid="53" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:21.00" />
                    <SPLIT distance="150" swimtime="00:02:05.57" />
                    <SPLIT distance="200" swimtime="00:02:51.38" />
                    <SPLIT distance="250" swimtime="00:03:37.66" />
                    <SPLIT distance="300" swimtime="00:04:24.04" />
                    <SPLIT distance="350" swimtime="00:05:09.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="12" points="239" swimtime="00:01:28.41" resultid="175810154" heatid="65" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="216" swimtime="00:03:17.98" resultid="175810155" heatid="72" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.31" />
                    <SPLIT distance="100" swimtime="00:01:34.87" />
                    <SPLIT distance="150" swimtime="00:02:26.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Gajdowska" birthdate="1995-05-14" gender="F" nation="POL" license="102001600173" swrid="4258728" athleteid="4258728">
              <RESULTS>
                <RESULT eventid="2" points="579" swimtime="00:00:27.51" resultid="175810177" heatid="15" lane="4" />
                <RESULT eventid="4" points="618" swimtime="00:00:58.97" resultid="175810179" heatid="23" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" points="601" swimtime="00:02:10.66" resultid="175810178" heatid="37" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                    <SPLIT distance="100" swimtime="00:01:03.09" />
                    <SPLIT distance="150" swimtime="00:01:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="557" swimtime="00:01:08.68" resultid="175810180" heatid="146" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Romuald" lastname="Kozłowski" birthdate="1966-08-13" gender="M" nation="POL" license="512914700012" swrid="5425564" athleteid="5425564">
              <RESULTS>
                <RESULT eventid="1" points="354" swimtime="00:00:28.49" resultid="175810181" heatid="12" lane="6" />
                <RESULT eventid="16" points="382" swimtime="00:00:34.36" resultid="175810182" heatid="84" lane="4" />
                <RESULT eventid="18" points="373" swimtime="00:01:16.73" resultid="175810183" heatid="95" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="331" swimtime="00:01:11.19" resultid="175810184" heatid="142" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" license="510414700009" swrid="4655152" athleteid="4655152">
              <RESULTS>
                <RESULT eventid="1" points="161" swimtime="00:00:37.00" resultid="175810189" heatid="19" lane="4" />
                <RESULT eventid="3" points="144" swimtime="00:01:25.45" resultid="175810191" heatid="29" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="93" swimtime="00:03:39.19" resultid="175810190" heatid="44" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.43" />
                    <SPLIT distance="100" swimtime="00:01:44.45" />
                    <SPLIT distance="150" swimtime="00:02:43.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="104" swimtime="00:01:44.61" resultid="175810192" heatid="139" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Piaściński" birthdate="1976-09-19" gender="M" nation="POL" swrid="5626929" athleteid="5626929">
              <RESULTS>
                <RESULT eventid="3" points="384" swimtime="00:01:01.68" resultid="175810171" heatid="20" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="365" swimtime="00:02:18.96" resultid="175810170" heatid="42" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:05.97" />
                    <SPLIT distance="150" swimtime="00:01:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11" points="366" swimtime="00:01:07.55" resultid="175810169" heatid="70" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="382" swimtime="00:01:07.91" resultid="175810172" heatid="147" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Kośmider" birthdate="1966-03-01" gender="M" nation="POL" license="512914700009" swrid="4992964" athleteid="4992964">
              <RESULTS>
                <RESULT eventid="5" points="302" swimtime="00:02:27.96" resultid="175810161" heatid="42" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                    <SPLIT distance="150" swimtime="00:01:51.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="293" swimtime="00:05:19.31" resultid="175810164" heatid="52" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:17.44" />
                    <SPLIT distance="150" swimtime="00:01:57.39" />
                    <SPLIT distance="200" swimtime="00:02:37.82" />
                    <SPLIT distance="250" swimtime="00:03:18.32" />
                    <SPLIT distance="300" swimtime="00:03:59.41" />
                    <SPLIT distance="350" swimtime="00:04:40.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="263" swimtime="00:03:07.47" resultid="175810162" heatid="110" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.12" />
                    <SPLIT distance="100" swimtime="00:01:30.29" />
                    <SPLIT distance="150" swimtime="00:02:17.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="25" points="138" swimtime="00:03:29.19" resultid="175810163" heatid="130" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                    <SPLIT distance="100" swimtime="00:01:41.75" />
                    <SPLIT distance="150" swimtime="00:02:38.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Korpetta" birthdate="1959-12-27" gender="M" nation="POL" license="112914700013" swrid="4754654" athleteid="4754654">
              <RESULTS>
                <RESULT eventid="5" points="180" swimtime="00:02:55.77" resultid="175810174" heatid="43" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:22.95" />
                    <SPLIT distance="150" swimtime="00:02:09.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="158" swimtime="00:06:32.56" resultid="175810176" heatid="47" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                    <SPLIT distance="100" swimtime="00:01:32.49" />
                    <SPLIT distance="150" swimtime="00:02:24.19" />
                    <SPLIT distance="200" swimtime="00:03:16.02" />
                    <SPLIT distance="250" swimtime="00:04:09.24" />
                    <SPLIT distance="300" swimtime="00:05:01.21" />
                    <SPLIT distance="350" swimtime="00:05:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11" points="144" swimtime="00:01:32.01" resultid="175810173" heatid="64" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="138" swimtime="00:03:23.99" resultid="175810175" heatid="73" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.11" />
                    <SPLIT distance="100" swimtime="00:01:39.23" />
                    <SPLIT distance="150" swimtime="00:02:33.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arkadiusz" lastname="Aptewicz" birthdate="1993-12-20" gender="M" nation="POL" license="507414700150" swrid="4806379" athleteid="4806379">
              <RESULTS>
                <RESULT eventid="7" points="595" swimtime="00:04:12.24" resultid="175810160" heatid="52" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                    <SPLIT distance="100" swimtime="00:00:59.07" />
                    <SPLIT distance="150" swimtime="00:01:31.27" />
                    <SPLIT distance="200" swimtime="00:02:03.45" />
                    <SPLIT distance="250" swimtime="00:02:35.94" />
                    <SPLIT distance="300" swimtime="00:03:08.44" />
                    <SPLIT distance="350" swimtime="00:03:40.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="545" swimtime="00:00:30.54" resultid="175810157" heatid="89" lane="2" />
                <RESULT eventid="18" points="591" swimtime="00:01:05.84" resultid="175810159" heatid="95" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="626" swimtime="00:02:20.44" resultid="175810158" heatid="105" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:07.42" />
                    <SPLIT distance="150" swimtime="00:01:43.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kaczmarek" birthdate="1977-06-25" gender="M" nation="POL" license="512914700003" swrid="4043251" athleteid="4043251">
              <RESULTS>
                <RESULT eventid="9" points="569" swimtime="00:00:26.81" resultid="175810168" heatid="59" lane="3" />
                <RESULT eventid="11" points="545" swimtime="00:00:59.16" resultid="175810165" heatid="70" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="583" swimtime="00:00:26.03" resultid="175810167" heatid="117" lane="3" />
                <RESULT eventid="24" points="545" swimtime="00:00:58.49" resultid="175810166" heatid="125" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Brozyna" birthdate="1980-04-28" gender="M" nation="POL" license="512914700006" swrid="5312396" athleteid="5312396">
              <RESULTS>
                <RESULT eventid="9" points="282" swimtime="00:00:33.86" resultid="175810196" heatid="59" lane="6" />
                <RESULT eventid="11" points="291" swimtime="00:01:12.86" resultid="175810193" heatid="70" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="307" swimtime="00:02:36.47" resultid="175810195" heatid="73" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:01:16.98" />
                    <SPLIT distance="150" swimtime="00:01:57.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" points="325" swimtime="00:02:39.45" resultid="175810194" heatid="136" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="150" swimtime="00:02:02.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Timea Beatrix" lastname="Balajcza" birthdate="1971-09-22" gender="F" nation="POL" license="510414600003" swrid="5240601" athleteid="5240601">
              <RESULTS>
                <RESULT eventid="15" points="396" swimtime="00:00:38.88" resultid="175810145" heatid="80" lane="3" />
                <RESULT eventid="17" points="358" swimtime="00:01:27.76" resultid="175810147" heatid="101" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="349" swimtime="00:03:11.11" resultid="175810146" heatid="112" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="100" swimtime="00:01:30.60" />
                    <SPLIT distance="150" swimtime="00:02:20.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="298" swimtime="00:01:24.60" resultid="175810148" heatid="138" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Szyszkowska" birthdate="1996-11-05" gender="F" nation="POL" swrid="4282341" athleteid="4282341">
              <RESULTS>
                <RESULT eventid="15" points="556" swimtime="00:00:34.72" resultid="175810185" heatid="88" lane="4" />
                <RESULT eventid="17" points="554" swimtime="00:01:15.91" resultid="175810187" heatid="101" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="547" swimtime="00:02:44.53" resultid="175810186" heatid="112" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:20.31" />
                    <SPLIT distance="150" swimtime="00:02:02.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="524" swimtime="00:01:10.06" resultid="175810188" heatid="146" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="31" points="613" swimtime="00:01:43.44" resultid="175810197" heatid="149" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                    <SPLIT distance="100" swimtime="00:00:54.78" />
                    <SPLIT distance="150" swimtime="00:01:19.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4282341" number="1" />
                    <RELAYPOSITION athleteid="4258728" number="2" />
                    <RELAYPOSITION athleteid="4043251" number="3" />
                    <RELAYPOSITION athleteid="4806379" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="31" points="427" swimtime="00:01:56.66" resultid="175810199" heatid="149" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                    <SPLIT distance="100" swimtime="00:00:59.51" />
                    <SPLIT distance="150" swimtime="00:01:28.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4251116" number="1" />
                    <RELAYPOSITION athleteid="5626929" number="2" />
                    <RELAYPOSITION athleteid="5240932" number="3" />
                    <RELAYPOSITION athleteid="5425564" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="585" swimtime="00:01:54.97" resultid="175810198" heatid="153" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                    <SPLIT distance="100" swimtime="00:00:57.64" />
                    <SPLIT distance="150" swimtime="00:01:27.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4043251" number="1" />
                    <RELAYPOSITION athleteid="4806379" number="2" />
                    <RELAYPOSITION athleteid="4282341" number="3" />
                    <RELAYPOSITION athleteid="4258728" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="369" swimtime="00:02:14.08" resultid="175810200" heatid="153" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:12.58" />
                    <SPLIT distance="150" swimtime="00:01:43.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5240932" number="1" />
                    <RELAYPOSITION athleteid="5240601" number="2" />
                    <RELAYPOSITION athleteid="5425564" number="3" />
                    <RELAYPOSITION athleteid="4992964" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01506" nation="POL" region="06" clubid="90256" swrid="90256" name="BOSiR Brzesko">
          <ATHLETES>
            <ATHLETE firstname="Przemysław" lastname="Jurek" birthdate="1981-04-11" gender="M" nation="POL" swrid="4992923" athleteid="4992923">
              <RESULTS>
                <RESULT eventid="3" points="393" swimtime="00:01:01.17" resultid="175810144" heatid="33" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="400" swimtime="00:00:29.50" resultid="175810143" heatid="117" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03706" nation="POL" region="06" clubid="87567" swrid="87567" name="Stow. Siemacha ASP Kraków" shortname="Siemacha ASP Kraków">
          <ATHLETES>
            <ATHLETE firstname="Paulina" lastname="Palmowska" birthdate="1985-08-01" gender="F" nation="POL" license="503706600141" swrid="4992815" athleteid="4992815">
              <RESULTS>
                <RESULT eventid="6" points="381" swimtime="00:02:32.07" resultid="175810492" heatid="45" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:01:12.85" />
                    <SPLIT distance="150" swimtime="00:01:52.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10" points="442" swimtime="00:00:33.17" resultid="175810494" heatid="58" lane="4" />
                <RESULT eventid="12" points="420" swimtime="00:01:13.25" resultid="175810491" heatid="65" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="412" swimtime="00:02:39.79" resultid="175810493" heatid="72" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:17.07" />
                    <SPLIT distance="150" swimtime="00:01:58.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06711" nation="POL" region="11" clubid="67997" swrid="67997" name="Uczniowski Klub Sportowy Dragon">
          <ATHLETES>
            <ATHLETE firstname="Emil" lastname="Strumiński" birthdate="1988-05-18" gender="M" nation="POL" license="306711700032" swrid="5448220" athleteid="5448220">
              <RESULTS>
                <RESULT eventid="3" points="523" swimtime="00:00:55.62" resultid="175810583" heatid="30" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="526" swimtime="00:02:03.10" resultid="175810581" heatid="39" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                    <SPLIT distance="100" swimtime="00:00:59.62" />
                    <SPLIT distance="150" swimtime="00:01:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="485" swimtime="00:04:30.00" resultid="175810584" heatid="46" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                    <SPLIT distance="100" swimtime="00:01:03.45" />
                    <SPLIT distance="150" swimtime="00:01:37.87" />
                    <SPLIT distance="200" swimtime="00:02:13.06" />
                    <SPLIT distance="250" swimtime="00:02:47.95" />
                    <SPLIT distance="300" swimtime="00:03:22.74" />
                    <SPLIT distance="350" swimtime="00:03:57.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" points="459" swimtime="00:01:01.91" resultid="175810582" heatid="125" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06306" nation="POL" region="06" clubid="93235" swrid="93235" name="KS Korona 1919 Kraków" shortname="Korona 1919 Kraków">
          <ATHLETES>
            <ATHLETE firstname="Adam" lastname="Pycia" birthdate="1966-02-21" gender="M" nation="POL" swrid="4992712" athleteid="4992712">
              <RESULTS>
                <RESULT eventid="1" points="257" swimtime="00:00:31.67" resultid="175809974" heatid="6" lane="5" />
                <RESULT eventid="3" points="264" swimtime="00:01:09.81" resultid="175809976" heatid="28" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="236" swimtime="00:00:40.34" resultid="175809975" heatid="83" lane="1" />
                <RESULT eventid="30" points="194" swimtime="00:01:24.99" resultid="175809977" heatid="139" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Baranik" birthdate="1969-06-29" gender="M" nation="POL" license="506306700027" swrid="4992740" athleteid="4992740">
              <RESULTS>
                <RESULT eventid="1" points="412" swimtime="00:00:27.08" resultid="175809978" heatid="12" lane="3" />
                <RESULT eventid="22" points="395" swimtime="00:00:29.63" resultid="175809980" heatid="120" lane="4" />
                <RESULT eventid="24" points="252" swimtime="00:01:15.59" resultid="175809979" heatid="126" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="312" swimtime="00:01:12.64" resultid="175809981" heatid="140" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Leńczowska" birthdate="1982-01-15" gender="F" nation="POL" swrid="4992907" athleteid="4992907">
              <RESULTS>
                <RESULT eventid="2" points="372" swimtime="00:00:31.88" resultid="175809983" heatid="4" lane="2" />
                <RESULT eventid="10" points="302" swimtime="00:00:37.64" resultid="175809986" heatid="58" lane="2" />
                <RESULT eventid="12" points="297" swimtime="00:01:22.22" resultid="175809984" heatid="65" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="302" swimtime="00:02:57.24" resultid="175809985" heatid="74" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                    <SPLIT distance="100" swimtime="00:01:26.44" />
                    <SPLIT distance="150" swimtime="00:02:12.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Próchniewicz" birthdate="1978-02-18" gender="M" nation="POL" swrid="4992816" athleteid="4992816">
              <RESULTS>
                <RESULT eventid="1" points="158" swimtime="00:00:37.28" resultid="175809991" heatid="13" lane="3" />
                <RESULT eventid="9" points="75" swimtime="00:00:52.60" resultid="175809993" heatid="60" lane="2" />
                <RESULT eventid="30" points="81" swimtime="00:01:53.53" resultid="175809992" heatid="140" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Mleczko" birthdate="1947-08-26" gender="M" nation="POL" swrid="4992812" athleteid="4992812">
              <RESULTS>
                <RESULT eventid="1" points="131" swimtime="00:00:39.67" resultid="175809994" heatid="14" lane="6" />
                <RESULT eventid="3" points="136" swimtime="00:01:27.19" resultid="175809996" heatid="29" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="94" swimtime="00:03:38.44" resultid="175809995" heatid="40" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.45" />
                    <SPLIT distance="100" swimtime="00:01:50.63" />
                    <SPLIT distance="150" swimtime="00:02:45.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="90" swimtime="00:07:51.91" resultid="175809997" heatid="46" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.28" />
                    <SPLIT distance="100" swimtime="00:01:50.28" />
                    <SPLIT distance="150" swimtime="00:02:49.39" />
                    <SPLIT distance="200" swimtime="00:03:49.33" />
                    <SPLIT distance="250" swimtime="00:04:51.65" />
                    <SPLIT distance="300" swimtime="00:05:52.35" />
                    <SPLIT distance="350" swimtime="00:06:54.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariola" lastname="Kuliś" birthdate="1966-07-27" gender="F" nation="POL" swrid="4992797" athleteid="4992797">
              <RESULTS>
                <RESULT eventid="2" points="394" swimtime="00:00:31.26" resultid="175810007" heatid="4" lane="4" />
                <RESULT eventid="15" points="423" swimtime="00:00:38.02" resultid="175810008" heatid="80" lane="4" />
                <RESULT eventid="21" points="370" swimtime="00:00:33.94" resultid="175810009" heatid="113" lane="6" />
                <RESULT eventid="29" points="376" swimtime="00:01:18.29" resultid="175810010" heatid="143" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Damian" lastname="Kaczor" birthdate="1994-04-11" gender="M" nation="POL" swrid="4180452" athleteid="4180452">
              <RESULTS>
                <RESULT eventid="1" points="525" swimtime="00:00:24.99" resultid="175810017" heatid="8" lane="2" />
                <RESULT eventid="3" points="562" swimtime="00:00:54.31" resultid="175810019" heatid="30" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="534" swimtime="00:00:30.74" resultid="175810018" heatid="84" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Łysiak" birthdate="1973-03-30" gender="M" nation="POL" swrid="5468085" athleteid="5468085">
              <RESULTS>
                <RESULT eventid="1" points="258" swimtime="00:00:31.64" resultid="175810020" heatid="6" lane="4" />
                <RESULT eventid="5" points="242" swimtime="00:02:39.33" resultid="175810021" heatid="36" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:17.83" />
                    <SPLIT distance="150" swimtime="00:01:59.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="204" swimtime="00:00:37.74" resultid="175810023" heatid="60" lane="5" />
                <RESULT eventid="22" points="221" swimtime="00:00:35.95" resultid="175810022" heatid="121" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogusław" lastname="Kwiatkowski" birthdate="1956-07-24" gender="M" nation="POL" swrid="5468084" athleteid="5468084">
              <RESULTS>
                <RESULT eventid="1" points="70" swimtime="00:00:48.86" resultid="175810024" heatid="14" lane="5" />
                <RESULT eventid="3" points="65" swimtime="00:01:51.24" resultid="175810026" heatid="31" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="65" swimtime="00:04:06.95" resultid="175810025" heatid="36" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.05" />
                    <SPLIT distance="100" swimtime="00:01:54.09" />
                    <SPLIT distance="150" swimtime="00:03:01.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="60" swimtime="00:09:01.63" resultid="175810027" heatid="50" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.83" />
                    <SPLIT distance="100" swimtime="00:02:03.92" />
                    <SPLIT distance="150" swimtime="00:03:16.39" />
                    <SPLIT distance="200" swimtime="00:04:26.14" />
                    <SPLIT distance="250" swimtime="00:05:36.56" />
                    <SPLIT distance="300" swimtime="00:06:44.08" />
                    <SPLIT distance="350" swimtime="00:07:51.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Macierzewska" birthdate="1960-04-20" gender="F" nation="POL" swrid="4992827" athleteid="4992827">
              <RESULTS>
                <RESULT eventid="4" points="257" swimtime="00:01:18.95" resultid="175809989" heatid="22" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" points="261" swimtime="00:02:52.58" resultid="175809987" heatid="38" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:22.88" />
                    <SPLIT distance="150" swimtime="00:02:08.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" points="212" swimtime="00:01:31.45" resultid="175809988" heatid="123" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="26" points="197" swimtime="00:03:25.50" resultid="175809990" heatid="129" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                    <SPLIT distance="100" swimtime="00:01:37.00" />
                    <SPLIT distance="150" swimtime="00:02:31.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Zadrożny" birthdate="1966-12-07" gender="M" nation="POL" swrid="4992825" athleteid="4992825">
              <RESULTS>
                <RESULT eventid="3" points="162" swimtime="00:01:22.12" resultid="175810005" heatid="21" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="158" swimtime="00:06:31.86" resultid="175810006" heatid="46" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                    <SPLIT distance="100" swimtime="00:01:31.80" />
                    <SPLIT distance="150" swimtime="00:02:20.84" />
                    <SPLIT distance="200" swimtime="00:03:10.55" />
                    <SPLIT distance="250" swimtime="00:04:01.96" />
                    <SPLIT distance="300" swimtime="00:04:53.31" />
                    <SPLIT distance="350" swimtime="00:05:44.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Malgorzata" lastname="Orlewicz-Musial" birthdate="1960-05-29" gender="F" nation="POL" swrid="5352178" athleteid="5352178">
              <RESULTS>
                <RESULT eventid="8" points="92" swimtime="00:08:37.87" resultid="175810031" heatid="51" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.06" />
                    <SPLIT distance="100" swimtime="00:01:59.30" />
                    <SPLIT distance="150" swimtime="00:03:03.78" />
                    <SPLIT distance="200" swimtime="00:04:09.19" />
                    <SPLIT distance="250" swimtime="00:05:15.01" />
                    <SPLIT distance="300" swimtime="00:06:22.65" />
                    <SPLIT distance="350" swimtime="00:07:29.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="12" points="58" swimtime="00:02:21.38" resultid="175810028" heatid="68" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="27" points="70" swimtime="00:04:54.76" resultid="175810029" heatid="134" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.05" />
                    <SPLIT distance="100" swimtime="00:02:22.89" />
                    <SPLIT distance="150" swimtime="00:03:50.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="72" swimtime="00:02:15.65" resultid="175810030" heatid="145" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Janeczko" birthdate="1972-12-23" gender="F" nation="POL" swrid="4218717" athleteid="4218717">
              <RESULTS>
                <RESULT eventid="10" points="242" swimtime="00:00:40.50" resultid="175810004" heatid="58" lane="6" />
                <RESULT eventid="12" points="188" swimtime="00:01:35.79" resultid="175810001" heatid="68" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" points="278" swimtime="00:00:37.33" resultid="175810003" heatid="116" lane="4" />
                <RESULT eventid="23" points="195" swimtime="00:01:34.03" resultid="175810002" heatid="123" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Jawień" birthdate="1971-06-11" gender="M" nation="POL" swrid="5468083" athleteid="5468083">
              <RESULTS>
                <RESULT eventid="11" points="265" swimtime="00:01:15.19" resultid="175809970" heatid="67" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="251" swimtime="00:02:47.31" resultid="175809973" heatid="73" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:21.83" />
                    <SPLIT distance="150" swimtime="00:02:05.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" points="337" swimtime="00:01:19.41" resultid="175809972" heatid="99" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="320" swimtime="00:02:55.66" resultid="175809971" heatid="107" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:25.57" />
                    <SPLIT distance="150" swimtime="00:02:10.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Mucha" birthdate="1967-04-24" gender="M" nation="POL" swrid="4218718" athleteid="4218718">
              <RESULTS>
                <RESULT eventid="16" points="276" swimtime="00:00:38.28" resultid="175809982" heatid="87" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Bielańska-Bugiel" birthdate="1984-04-20" gender="F" nation="POL" swrid="5468078" athleteid="5468078">
              <RESULTS>
                <RESULT eventid="15" points="110" swimtime="00:00:59.60" resultid="175810011" heatid="86" lane="6" />
                <RESULT eventid="19" points="110" swimtime="00:04:40.07" resultid="175810012" heatid="108" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.60" />
                    <SPLIT distance="100" swimtime="00:02:13.42" />
                    <SPLIT distance="150" swimtime="00:03:29.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Toporski" birthdate="1959-10-20" gender="M" nation="POL" swrid="5484421" athleteid="5484421">
              <RESULTS>
                <RESULT eventid="18" points="147" swimtime="00:01:44.56" resultid="175810015" heatid="100" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="163" swimtime="00:03:39.57" resultid="175810014" heatid="103" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.91" />
                    <SPLIT distance="100" swimtime="00:01:47.15" />
                    <SPLIT distance="150" swimtime="00:02:44.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" points="75" swimtime="00:01:53.11" resultid="175810013" heatid="127" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="25" points="81" swimtime="00:04:09.53" resultid="175810016" heatid="130" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.16" />
                    <SPLIT distance="100" swimtime="00:02:00.11" />
                    <SPLIT distance="150" swimtime="00:03:06.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Romańska" birthdate="1975-04-22" gender="F" nation="POL" swrid="4992818" athleteid="4992818">
              <RESULTS>
                <RESULT eventid="21" points="85" swimtime="00:00:55.40" resultid="175809999" heatid="116" lane="5" />
                <RESULT eventid="27" points="116" swimtime="00:04:09.82" resultid="175809998" heatid="134" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.70" />
                    <SPLIT distance="100" swimtime="00:02:06.42" />
                    <SPLIT distance="150" swimtime="00:03:14.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="117" swimtime="00:01:55.38" resultid="175810000" heatid="145" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="31" points="302" swimtime="00:02:10.94" resultid="175810032" heatid="148" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:05.44" />
                    <SPLIT distance="150" swimtime="00:01:32.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4992797" number="1" />
                    <RELAYPOSITION athleteid="4992827" number="2" />
                    <RELAYPOSITION athleteid="4992740" number="3" />
                    <RELAYPOSITION athleteid="4992812" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="31" points="108" swimtime="00:03:04.16" resultid="175810034" heatid="150" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.15" />
                    <SPLIT distance="100" swimtime="00:01:32.71" />
                    <SPLIT distance="150" swimtime="00:02:22.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5468084" number="1" />
                    <RELAYPOSITION athleteid="4992818" number="2" />
                    <RELAYPOSITION athleteid="5352178" number="3" />
                    <RELAYPOSITION athleteid="5484421" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="31" points="296" swimtime="00:02:11.79" resultid="175810036" heatid="150" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:02.93" />
                    <SPLIT distance="150" swimtime="00:01:37.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4992907" number="1" />
                    <RELAYPOSITION athleteid="5468083" number="2" />
                    <RELAYPOSITION athleteid="4218717" number="3" />
                    <RELAYPOSITION athleteid="4218718" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="128" swimtime="00:03:10.71" resultid="175810033" heatid="151" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                    <SPLIT distance="100" swimtime="00:01:30.82" />
                    <SPLIT distance="150" swimtime="00:02:24.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4992827" number="1" />
                    <RELAYPOSITION athleteid="5484421" number="2" />
                    <RELAYPOSITION athleteid="4992818" number="3" />
                    <RELAYPOSITION athleteid="5468084" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" points="354" swimtime="00:02:15.88" resultid="175810035" heatid="152" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:01:14.66" />
                    <SPLIT distance="150" swimtime="00:01:44.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4992907" number="1" />
                    <RELAYPOSITION athleteid="5468083" number="2" />
                    <RELAYPOSITION athleteid="4992740" number="3" />
                    <RELAYPOSITION athleteid="4992797" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02202" nation="POL" region="02" clubid="87558" swrid="87558" name="MKS Astoria Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-13" gender="M" nation="POL" license="102202700126" swrid="5471726" athleteid="5471726">
              <RESULTS>
                <RESULT eventid="9" points="89" swimtime="00:00:49.71" resultid="175809859" heatid="56" lane="2" />
                <RESULT eventid="11" points="86" swimtime="00:01:49.09" resultid="175809856" heatid="63" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="74" swimtime="00:04:10.90" resultid="175809858" heatid="71" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.20" />
                    <SPLIT distance="100" swimtime="00:02:00.81" />
                    <SPLIT distance="150" swimtime="00:03:04.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" points="156" swimtime="00:00:46.30" resultid="175809857" heatid="79" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08114" nation="POL" region="14" clubid="90775" swrid="90775" name="KU AZS Uniwersytetu Warszawskiego" name.en="Ku Azs Uw">
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Rębas" birthdate="1989-12-11" gender="M" nation="POL" license="508114700069" swrid="4251117" athleteid="4251117">
              <RESULTS>
                <RESULT eventid="1" points="487" swimtime="00:00:25.61" resultid="175810460" heatid="8" lane="3" />
                <RESULT eventid="3" points="539" swimtime="00:00:55.07" resultid="175810462" heatid="30" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" points="504" swimtime="00:01:00.03" resultid="175810461" heatid="125" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="25" points="477" swimtime="00:02:18.50" resultid="175810463" heatid="130" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                    <SPLIT distance="100" swimtime="00:01:04.79" />
                    <SPLIT distance="150" swimtime="00:01:40.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02801" nation="POL" region="01" clubid="85848" swrid="85848" name="KS Masters Polkowice" shortname="Masters Polkowice">
          <ATHLETES>
            <ATHLETE firstname="Pavlo" lastname="Vechirko" birthdate="1968-01-02" gender="M" nation="POL" swrid="5626940" athleteid="5626940">
              <RESULTS>
                <RESULT eventid="9" points="225" swimtime="00:00:36.50" resultid="175810106" heatid="55" lane="5" />
                <RESULT eventid="11" points="237" swimtime="00:01:18.03" resultid="175810103" heatid="67" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" points="274" swimtime="00:01:25.02" resultid="175810105" heatid="96" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="260" swimtime="00:03:08.04" resultid="175810104" heatid="110" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                    <SPLIT distance="100" swimtime="00:01:30.88" />
                    <SPLIT distance="150" swimtime="00:02:19.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" region="11" clubid="65759" swrid="65759" name="KS Górnik Radlin">
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Kubica" birthdate="1972-02-22" gender="M" nation="POL" swrid="5398297" athleteid="5398297">
              <RESULTS>
                <RESULT eventid="11" points="249" swimtime="00:01:16.82" resultid="175810212" heatid="67" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="303" swimtime="00:00:32.35" resultid="175810214" heatid="114" lane="4" />
                <RESULT eventid="24" points="274" swimtime="00:01:13.52" resultid="175810213" heatid="126" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="25" points="227" swimtime="00:02:57.30" resultid="175810215" heatid="128" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                    <SPLIT distance="100" swimtime="00:01:21.66" />
                    <SPLIT distance="150" swimtime="00:02:09.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01911" nation="POL" region="11" clubid="67927" swrid="67927" name="RMKS Rybnik">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Duda" birthdate="1981-04-15" gender="F" nation="POL" swrid="4992966" athleteid="4992966">
              <RESULTS>
                <RESULT eventid="2" points="477" swimtime="00:00:29.34" resultid="175810201" heatid="15" lane="1" />
                <RESULT eventid="4" points="428" swimtime="00:01:06.65" resultid="175810204" heatid="23" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" points="371" swimtime="00:00:39.72" resultid="175810202" heatid="80" lane="1" />
                <RESULT eventid="21" points="430" swimtime="00:00:32.29" resultid="175810203" heatid="113" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Henzel" birthdate="1971-09-20" gender="M" nation="POL" swrid="5626907" athleteid="5626907">
              <RESULTS>
                <RESULT eventid="3" points="179" swimtime="00:01:19.51" resultid="175810206" heatid="25" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="127" swimtime="00:00:43.18" resultid="175810205" heatid="122" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Rodak" birthdate="1982-08-02" gender="M" nation="POL" swrid="5626932" athleteid="5626932">
              <RESULTS>
                <RESULT eventid="3" points="93" swimtime="00:01:38.62" resultid="175810207" heatid="32" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marlena" lastname="Stephan" birthdate="1975-02-20" gender="F" nation="POL" swrid="5626936" athleteid="5626936">
              <RESULTS>
                <RESULT eventid="15" points="166" swimtime="00:00:51.87" resultid="175810208" heatid="77" lane="2" />
                <RESULT eventid="17" points="140" swimtime="00:02:00.02" resultid="175810209" heatid="91" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="126" swimtime="00:01:52.47" resultid="175810210" heatid="145" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="32" points="174" swimtime="00:02:52.14" resultid="175810211" heatid="151" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4992966" number="1" />
                    <RELAYPOSITION athleteid="5626907" number="2" />
                    <RELAYPOSITION athleteid="5626932" number="3" />
                    <RELAYPOSITION athleteid="5626936" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="07611" nation="POL" region="11" clubid="77420" swrid="77420" name="Uks Dragon">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Jankowski" birthdate="1995-08-14" gender="M" nation="POL" swrid="4112623" athleteid="4112623">
              <RESULTS>
                <RESULT eventid="3" points="664" swimtime="00:00:51.38" resultid="175810097" heatid="30" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="656" swimtime="00:00:25.56" resultid="175810098" heatid="59" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00201" nation="POL" region="01" clubid="65762" swrid="65762" name="KS AZS AWF Wrocław" shortname="AZS AWF Wroclaw">
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Sasin" birthdate="1994-04-15" gender="F" nation="POL" license="100201600097" swrid="4236079" athleteid="4236079">
              <RESULTS>
                <RESULT eventid="6" points="570" swimtime="00:02:13.01" resultid="175809860" heatid="37" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:03.41" />
                    <SPLIT distance="150" swimtime="00:01:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" points="588" swimtime="00:01:05.13" resultid="175809861" heatid="123" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01610" nation="POL" region="10" clubid="75878" swrid="75878" name="Grupa Pływacka Gdynia Masters" shortname="Masters Gdynia">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Gorbaczow" birthdate="1958-12-28" gender="M" nation="POL" swrid="4191113" athleteid="4191113">
              <RESULTS>
                <RESULT eventid="1" points="296" swimtime="00:00:30.25" resultid="175809836" heatid="2" lane="6" />
                <RESULT eventid="3" points="306" swimtime="00:01:06.49" resultid="175809838" heatid="20" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="283" swimtime="00:02:31.23" resultid="175809837" heatid="35" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:14.27" />
                    <SPLIT distance="150" swimtime="00:01:53.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="258" swimtime="00:00:34.89" resultid="175809839" heatid="55" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05911" nation="POL" region="11" clubid="89648" swrid="89648" name="UKS Karlik Katowice">
          <ATHLETES>
            <ATHLETE firstname="Karolina" lastname="Nowak" birthdate="1997-09-07" gender="F" nation="POL" swrid="5626927" athleteid="5626927">
              <RESULTS>
                <RESULT eventid="2" points="219" swimtime="00:00:38.01" resultid="175810385" heatid="9" lane="2" />
                <RESULT eventid="4" points="193" swimtime="00:01:26.95" resultid="175810387" heatid="22" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10" points="146" swimtime="00:00:47.90" resultid="175810388" heatid="61" lane="3" />
                <RESULT eventid="15" points="188" swimtime="00:00:49.82" resultid="175810386" heatid="85" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szczypiński" birthdate="1986-12-05" gender="M" nation="POL" swrid="4060998" athleteid="4060998">
              <RESULTS>
                <RESULT eventid="3" points="481" swimtime="00:00:57.22" resultid="175810383" heatid="33" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="466" swimtime="00:02:08.13" resultid="175810381" heatid="39" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:01.43" />
                    <SPLIT distance="150" swimtime="00:01:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="412" swimtime="00:00:29.86" resultid="175810384" heatid="55" lane="4" />
                <RESULT eventid="24" points="417" swimtime="00:01:03.93" resultid="175810382" heatid="126" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02611" nation="POL" region="11" clubid="74354" swrid="74354" name="Towarzystwo Sportowe Weteran Zabrze" shortname="TS Weteran Zabrze">
          <ATHLETES>
            <ATHLETE firstname="Wieslaw" lastname="Kornicki" birthdate="1949-01-28" gender="M" nation="POL" swrid="4137183" athleteid="4137183">
              <RESULTS>
                <RESULT eventid="1" points="177" swimtime="00:00:35.89" resultid="175810361" heatid="6" lane="6" />
                <RESULT eventid="16" points="128" swimtime="00:00:49.39" resultid="175810362" heatid="79" lane="6" />
                <RESULT eventid="22" points="170" swimtime="00:00:39.22" resultid="175810363" heatid="119" lane="2" />
                <RESULT eventid="30" points="119" swimtime="00:01:40.11" resultid="175810364" heatid="141" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Genowefa" lastname="Drużyńska" birthdate="1951-02-18" gender="F" nation="POL" swrid="4655173" athleteid="4655173">
              <RESULTS>
                <RESULT eventid="2" points="75" swimtime="00:00:54.33" resultid="175810365" heatid="16" lane="5" />
                <RESULT eventid="15" points="78" swimtime="00:01:06.81" resultid="175810366" heatid="78" lane="3" />
                <RESULT eventid="17" points="66" swimtime="00:02:33.76" resultid="175810367" heatid="91" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="69" swimtime="00:02:17.45" resultid="175810368" heatid="143" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wjciech" lastname="Kosiak" birthdate="1940-04-20" gender="M" nation="POL" swrid="5582455" athleteid="5582455">
              <RESULTS>
                <RESULT eventid="1" points="72" swimtime="00:00:48.25" resultid="175810377" heatid="14" lane="2" />
                <RESULT eventid="3" points="73" swimtime="00:01:46.91" resultid="175810380" heatid="31" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="63" swimtime="00:04:08.97" resultid="175810378" heatid="40" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.18" />
                    <SPLIT distance="100" swimtime="00:02:04.33" />
                    <SPLIT distance="150" swimtime="00:03:10.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="33" swimtime="00:01:07.70" resultid="175810379" heatid="115" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beata" lastname="Sulewska" birthdate="1972-11-02" gender="F" nation="POL" swrid="4792005" athleteid="4792005">
              <RESULTS>
                <RESULT eventid="6" points="421" swimtime="00:02:27.09" resultid="175810358" heatid="45" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:50.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8" points="432" swimtime="00:05:09.23" resultid="175810360" heatid="53" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:14.32" />
                    <SPLIT distance="150" swimtime="00:01:53.10" />
                    <SPLIT distance="200" swimtime="00:02:32.73" />
                    <SPLIT distance="250" swimtime="00:03:12.40" />
                    <SPLIT distance="300" swimtime="00:03:52.06" />
                    <SPLIT distance="350" swimtime="00:04:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="17" points="412" swimtime="00:01:23.78" resultid="175810359" heatid="101" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Twardysko" birthdate="1956-01-16" gender="M" nation="POL" swrid="5464152" athleteid="5464152">
              <RESULTS>
                <RESULT eventid="5" points="181" swimtime="00:02:55.41" resultid="175810370" heatid="43" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:01:23.68" />
                    <SPLIT distance="150" swimtime="00:02:09.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" points="166" swimtime="00:06:25.82" resultid="175810372" heatid="47" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:01:28.22" />
                    <SPLIT distance="150" swimtime="00:02:17.04" />
                    <SPLIT distance="200" swimtime="00:03:06.64" />
                    <SPLIT distance="250" swimtime="00:03:57.32" />
                    <SPLIT distance="300" swimtime="00:04:47.68" />
                    <SPLIT distance="350" swimtime="00:05:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11" points="132" swimtime="00:01:34.87" resultid="175810369" heatid="64" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="117" swimtime="00:03:35.74" resultid="175810371" heatid="71" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.64" />
                    <SPLIT distance="100" swimtime="00:01:42.62" />
                    <SPLIT distance="150" swimtime="00:02:40.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teresa" lastname="Żylińska" birthdate="1950-10-13" gender="F" nation="POL" swrid="5464154" athleteid="5464154">
              <RESULTS>
                <RESULT eventid="6" points="64" swimtime="00:04:35.39" resultid="175810374" heatid="41" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.00" />
                    <SPLIT distance="100" swimtime="00:02:11.75" />
                    <SPLIT distance="150" swimtime="00:03:25.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8" points="67" swimtime="00:09:35.50" resultid="175810376" heatid="49" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.64" />
                    <SPLIT distance="100" swimtime="00:02:12.58" />
                    <SPLIT distance="150" swimtime="00:03:27.23" />
                    <SPLIT distance="200" swimtime="00:04:41.25" />
                    <SPLIT distance="250" swimtime="00:05:55.29" />
                    <SPLIT distance="300" swimtime="00:07:10.03" />
                    <SPLIT distance="350" swimtime="00:08:23.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="12" points="64" swimtime="00:02:17.05" resultid="175810373" heatid="69" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="66" swimtime="00:04:53.68" resultid="175810375" heatid="74" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.81" />
                    <SPLIT distance="100" swimtime="00:02:23.16" />
                    <SPLIT distance="150" swimtime="00:03:40.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="65774" swrid="65774" name="KS WARTA Poznań">
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Lesinski" birthdate="1944-04-13" gender="M" nation="POL" swrid="4188190" athleteid="4188190">
              <RESULTS>
                <RESULT eventid="1" points="99" swimtime="00:00:43.49" resultid="175810445" heatid="14" lane="3" />
                <RESULT eventid="3" points="90" swimtime="00:01:39.82" resultid="175810447" heatid="31" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="93" swimtime="00:00:48.92" resultid="175810448" heatid="56" lane="5" />
                <RESULT eventid="11" points="83" swimtime="00:01:50.37" resultid="175810446" heatid="63" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Krupińska" birthdate="1953-05-24" gender="F" nation="POL" swrid="4992790" athleteid="4992790">
              <RESULTS>
                <RESULT eventid="4" points="64" swimtime="00:02:05.32" resultid="175810432" heatid="26" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" points="140" swimtime="00:00:55.00" resultid="175810430" heatid="86" lane="3" />
                <RESULT eventid="17" points="122" swimtime="00:02:05.45" resultid="175810433" heatid="98" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="130" swimtime="00:04:25.21" resultid="175810431" heatid="108" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.86" />
                    <SPLIT distance="100" swimtime="00:02:09.92" />
                    <SPLIT distance="150" swimtime="00:03:19.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Kotecka" birthdate="1965-05-08" gender="F" nation="POL" license="100115600357" swrid="4754727" athleteid="4754727">
              <RESULTS>
                <RESULT eventid="6" points="211" swimtime="00:03:05.00" resultid="175810438" heatid="45" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                    <SPLIT distance="100" swimtime="00:01:29.02" />
                    <SPLIT distance="150" swimtime="00:02:17.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8" points="220" swimtime="00:06:27.36" resultid="175810440" heatid="49" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                    <SPLIT distance="100" swimtime="00:01:30.32" />
                    <SPLIT distance="150" swimtime="00:02:19.21" />
                    <SPLIT distance="200" swimtime="00:03:08.98" />
                    <SPLIT distance="250" swimtime="00:03:59.74" />
                    <SPLIT distance="300" swimtime="00:04:49.69" />
                    <SPLIT distance="350" swimtime="00:05:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="12" points="159" swimtime="00:01:41.26" resultid="175810437" heatid="69" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="159" swimtime="00:03:39.30" resultid="175810439" heatid="72" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.02" />
                    <SPLIT distance="100" swimtime="00:01:47.76" />
                    <SPLIT distance="150" swimtime="00:02:43.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Szala" birthdate="1959-03-19" gender="F" nation="POL" swrid="4302573" athleteid="4302573">
              <RESULTS>
                <RESULT eventid="8" points="262" swimtime="00:06:05.48" resultid="175810443" heatid="53" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:27.54" />
                    <SPLIT distance="150" swimtime="00:02:14.15" />
                    <SPLIT distance="200" swimtime="00:03:00.85" />
                    <SPLIT distance="250" swimtime="00:03:47.46" />
                    <SPLIT distance="300" swimtime="00:04:33.87" />
                    <SPLIT distance="350" swimtime="00:05:20.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="12" points="234" swimtime="00:01:28.97" resultid="175810441" heatid="65" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="249" swimtime="00:03:08.83" resultid="175810442" heatid="72" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                    <SPLIT distance="100" swimtime="00:01:33.47" />
                    <SPLIT distance="150" swimtime="00:02:22.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="27" points="259" swimtime="00:03:11.00" resultid="175810444" heatid="135" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:31.03" />
                    <SPLIT distance="150" swimtime="00:02:25.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Waraczewski" birthdate="1962-04-19" gender="M" nation="POL" swrid="4992781" athleteid="4992781">
              <RESULTS>
                <RESULT eventid="16" points="254" swimtime="00:00:39.39" resultid="175810427" heatid="83" lane="4" />
                <RESULT eventid="18" points="254" swimtime="00:01:27.24" resultid="175810429" heatid="99" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="251" swimtime="00:03:10.43" resultid="175810428" heatid="107" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                    <SPLIT distance="100" swimtime="00:01:30.60" />
                    <SPLIT distance="150" swimtime="00:02:19.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystian" lastname="Talar" birthdate="2002-10-03" gender="M" nation="POL" swrid="4790712" athleteid="4790712">
              <RESULTS>
                <RESULT eventid="16" points="139" swimtime="00:00:48.11" resultid="175810434" heatid="84" lane="6" />
                <RESULT eventid="18" points="118" swimtime="00:01:52.40" resultid="175810436" heatid="96" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" points="114" swimtime="00:04:07.41" resultid="175810435" heatid="110" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.72" />
                    <SPLIT distance="100" swimtime="00:01:52.53" />
                    <SPLIT distance="150" swimtime="00:02:59.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Skurczyńska" birthdate="1971-10-13" gender="F" nation="POL" swrid="5626935" athleteid="5626935">
              <RESULTS>
                <RESULT eventid="15" points="210" swimtime="00:00:48.03" resultid="175810449" heatid="85" lane="2" />
                <RESULT eventid="19" points="174" swimtime="00:04:00.87" resultid="175810450" heatid="109" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.57" />
                    <SPLIT distance="100" swimtime="00:01:51.86" />
                    <SPLIT distance="150" swimtime="00:02:55.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="15" clubid="86433" swrid="86433" name="KU AZS U.A.M. Poznań">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Juszkiewicz" birthdate="1974-05-10" gender="M" nation="POL" license="503315700077" swrid="5537971" athleteid="5537971">
              <RESULTS>
                <RESULT eventid="1" points="265" swimtime="00:00:31.37" resultid="175810458" heatid="2" lane="1" />
                <RESULT eventid="5" points="232" swimtime="00:02:41.53" resultid="175810459" heatid="36" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="150" swimtime="00:02:02.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05806" nation="POL" region="06" clubid="93187" swrid="93187" name="IKS Druga Strona Sportu">
          <ATHLETES>
            <ATHLETE firstname="Tadeusz" lastname="Krawczyk" birthdate="1943-05-16" gender="M" nation="POL" swrid="4992809" athleteid="4992809">
              <RESULTS>
                <RESULT eventid="1" points="24" swimtime="00:01:09.89" resultid="175810599" heatid="14" lane="4" />
                <RESULT eventid="3" points="20" swimtime="00:02:45.04" resultid="175810601" heatid="29" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="18" swimtime="00:06:12.70" resultid="175810600" heatid="40" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.83" />
                    <SPLIT distance="100" swimtime="00:03:00.23" />
                    <SPLIT distance="150" swimtime="00:04:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9" points="14" swimtime="00:01:30.46" resultid="175810602" heatid="60" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogdan" lastname="Szczurek" birthdate="1952-02-07" gender="M" nation="POL" swrid="5626937" athleteid="5626937">
              <RESULTS>
                <RESULT eventid="3" points="60" swimtime="00:01:54.10" resultid="175810605" heatid="32" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="55" swimtime="00:04:21.21" resultid="175810604" heatid="36" lane="6" />
                <RESULT eventid="11" points="58" swimtime="00:02:04.16" resultid="175810603" heatid="66" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="62" swimtime="00:04:26.52" resultid="175810606" heatid="75" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.73" />
                    <SPLIT distance="100" swimtime="00:02:09.35" />
                    <SPLIT distance="150" swimtime="00:03:20.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Rupp" birthdate="1956-03-06" gender="F" nation="POL" swrid="5484417" athleteid="5484417">
              <RESULTS>
                <RESULT eventid="8" points="85" swimtime="00:08:50.51" resultid="175810598" heatid="49" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.62" />
                    <SPLIT distance="100" swimtime="00:02:02.58" />
                    <SPLIT distance="150" swimtime="00:03:11.42" />
                    <SPLIT distance="200" swimtime="00:04:18.55" />
                    <SPLIT distance="250" swimtime="00:05:25.93" />
                    <SPLIT distance="300" swimtime="00:06:34.70" />
                    <SPLIT distance="350" swimtime="00:07:42.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="12" points="65" swimtime="00:02:15.98" resultid="175810595" heatid="69" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" points="74" swimtime="00:04:42.23" resultid="175810597" heatid="74" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.71" />
                    <SPLIT distance="100" swimtime="00:02:15.77" />
                    <SPLIT distance="150" swimtime="00:03:30.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="27" points="68" swimtime="00:04:57.95" resultid="175810596" heatid="135" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.32" />
                    <SPLIT distance="100" swimtime="00:02:29.53" />
                    <SPLIT distance="150" swimtime="00:03:53.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00607" nation="POL" region="07" clubid="75298" swrid="75298" name="TP Masters Opole">
          <ATHLETES>
            <ATHLETE firstname="Jerzy" lastname="Minkiewicz" birthdate="1956-05-31" gender="M" nation="POL" swrid="4183581" athleteid="4183581">
              <RESULTS>
                <RESULT eventid="1" points="205" swimtime="00:00:34.18" resultid="175810351" heatid="11" lane="3" />
                <RESULT eventid="9" points="124" swimtime="00:00:44.46" resultid="175810353" heatid="57" lane="2" />
                <RESULT eventid="22" points="158" swimtime="00:00:40.20" resultid="175810352" heatid="119" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Mandziuk" birthdate="1965-04-11" gender="M" nation="POL" swrid="5626918" athleteid="5626918">
              <RESULTS>
                <RESULT eventid="1" points="178" swimtime="00:00:35.83" resultid="175810354" heatid="19" lane="3" />
                <RESULT eventid="3" points="168" swimtime="00:01:21.19" resultid="175810356" heatid="29" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="137" swimtime="00:03:12.43" resultid="175810355" heatid="43" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:01:29.11" />
                    <SPLIT distance="150" swimtime="00:02:22.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" points="104" status="DSQ" swimtime="00:01:57.36" resultid="175810357" heatid="100" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="14814" nation="POL" region="14" clubid="93424" swrid="93424" name="SP Legia Warszawa" shortname="Legia Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Grzelak" birthdate="1970-05-05" gender="M" nation="POL" swrid="4951293" athleteid="4951293">
              <RESULTS>
                <RESULT eventid="1" points="226" swimtime="00:00:33.07" resultid="175810099" heatid="3" lane="1" />
                <RESULT eventid="5" points="218" swimtime="00:02:45.06" resultid="175810100" heatid="40" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:20.62" />
                    <SPLIT distance="150" swimtime="00:02:03.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" points="217" swimtime="00:00:36.14" resultid="175810101" heatid="121" lane="4" />
                <RESULT eventid="25" points="159" swimtime="00:03:19.38" resultid="175810102" heatid="130" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                    <SPLIT distance="100" swimtime="00:01:32.60" />
                    <SPLIT distance="150" swimtime="00:02:26.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02706" nation="POL" region="06" clubid="82159" swrid="82159" name="UKS Jasień Sucha Beskidzka">
          <ATHLETES>
            <ATHLETE firstname="Aneta" lastname="Pytel" birthdate="1979-02-03" gender="F" nation="POL" swrid="5582461" athleteid="5582461">
              <RESULTS>
                <RESULT eventid="10" points="133" swimtime="00:00:49.44" resultid="175810590" heatid="61" lane="4" />
                <RESULT eventid="17" points="168" swimtime="00:01:52.82" resultid="175810589" heatid="98" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sabina" lastname="Sikora" birthdate="1984-10-03" gender="F" nation="POL" license="102706600159" swrid="5468086" athleteid="5468086">
              <RESULTS>
                <RESULT eventid="15" points="531" swimtime="00:00:35.26" resultid="175810591" heatid="88" lane="5" />
                <RESULT eventid="17" points="449" swimtime="00:01:21.43" resultid="175810593" heatid="101" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" points="375" swimtime="00:03:06.52" resultid="175810592" heatid="112" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                    <SPLIT distance="150" swimtime="00:02:19.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" points="426" swimtime="00:01:15.10" resultid="175810594" heatid="138" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00309" nation="POL" region="09" clubid="65783" swrid="65783" name="MKS JUVENIA Białystok">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Zmiejko" birthdate="1963-01-16" gender="M" nation="POL" swrid="4186249" athleteid="4186249">
              <RESULTS>
                <RESULT eventid="1" points="351" swimtime="00:00:28.57" resultid="175810454" heatid="17" lane="4" />
                <RESULT eventid="3" points="357" swimtime="00:01:03.18" resultid="175810456" heatid="34" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" points="321" swimtime="00:01:09.76" resultid="175810455" heatid="126" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="326" swimtime="00:01:11.58" resultid="175810457" heatid="147" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Michalik" birthdate="1979-07-14" gender="F" nation="POL" license="500309600228" swrid="4595750" athleteid="4595750">
              <RESULTS>
                <RESULT eventid="4" points="439" swimtime="00:01:06.09" resultid="175810452" heatid="23" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" points="460" swimtime="00:02:22.87" resultid="175810451" heatid="37" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                    <SPLIT distance="150" swimtime="00:01:45.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8" points="441" swimtime="00:05:07.19" resultid="175810453" heatid="53" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:14.41" />
                    <SPLIT distance="150" swimtime="00:01:53.52" />
                    <SPLIT distance="200" swimtime="00:02:32.58" />
                    <SPLIT distance="250" swimtime="00:03:11.91" />
                    <SPLIT distance="300" swimtime="00:03:50.74" />
                    <SPLIT distance="350" swimtime="00:04:29.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="07311" nation="POL" region="11" clubid="77475" swrid="77475" name="UKS &quot;Dwójeczka&quot; Częstochowa">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Lewiński" birthdate="1982-08-03" gender="M" nation="POL" swrid="5626915" athleteid="5626915">
              <RESULTS>
                <RESULT eventid="1" points="227" swimtime="00:00:33.02" resultid="175810093" heatid="13" lane="5" />
                <RESULT eventid="3" points="194" swimtime="00:01:17.34" resultid="175810095" heatid="32" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" points="161" swimtime="00:03:02.54" resultid="175810094" heatid="36" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                    <SPLIT distance="100" swimtime="00:01:21.84" />
                    <SPLIT distance="150" swimtime="00:02:12.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" points="175" swimtime="00:01:28.01" resultid="175810096" heatid="139" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ireneusz" lastname="Stachurski" birthdate="1969-07-22" gender="M" nation="POL" swrid="5464094" athleteid="5464094">
              <RESULTS>
                <RESULT eventid="7" points="185" swimtime="00:06:12.08" resultid="175810092" heatid="47" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="100" swimtime="00:01:25.89" />
                    <SPLIT distance="150" swimtime="00:02:14.62" />
                    <SPLIT distance="200" swimtime="00:03:03.52" />
                    <SPLIT distance="250" swimtime="00:03:51.67" />
                    <SPLIT distance="300" swimtime="00:04:40.16" />
                    <SPLIT distance="350" swimtime="00:05:28.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11" points="131" swimtime="00:01:34.97" resultid="175810089" heatid="63" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" points="134" swimtime="00:03:26.40" resultid="175810091" heatid="75" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.50" />
                    <SPLIT distance="100" swimtime="00:01:40.15" />
                    <SPLIT distance="150" swimtime="00:02:34.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" points="99" swimtime="00:01:43.20" resultid="175810090" heatid="124" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Michał Derewecki" version="11.69132">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Poznań" name="Letnie Mistrzostwa Okręgu Wielkopolskiego, Letnie Otwarte Korespondencyjne Mistrzostwa Polski w kategoriach Masters" course="LCM" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2021-06-26" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Poznań" nation="POL" />
      <POINTTABLE pointtableid="3014" name="FINA Point Scoring" version="2021" />
      <QUALIFY from="2020-03-01" until="2021-06-25" />
      <SESSIONS>
        <SESSION date="2021-06-26" daytime="09:15" endtime="16:09" number="1">
          <EVENTS>
            <EVENT eventid="1059" daytime="09:16" gender="X" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1060" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1885" />
                    <RANKING order="2" place="2" resultid="1883" />
                    <RANKING order="3" place="3" resultid="2356" />
                    <RANKING order="4" place="4" resultid="2184" />
                    <RANKING order="5" place="5" resultid="1599" />
                    <RANKING order="6" place="6" resultid="2357" />
                    <RANKING order="7" place="7" resultid="2185" />
                    <RANKING order="8" place="8" resultid="2358" />
                    <RANKING order="9" place="9" resultid="1884" />
                    <RANKING order="10" place="10" resultid="2094" />
                    <RANKING order="11" place="11" resultid="1600" />
                    <RANKING order="12" place="12" resultid="2355" />
                    <RANKING order="13" place="13" resultid="1958" />
                    <RANKING order="14" place="13" resultid="2095" />
                    <RANKING order="15" place="15" resultid="1251" />
                    <RANKING order="16" place="-1" resultid="1379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1061" agemax="16" agemin="14" />
                <AGEGROUP agegroupid="1062" agemax="13" agemin="10" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2947" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2948" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1063" daytime="09:20" gender="F" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2237" />
                    <RANKING order="2" place="2" resultid="2232" />
                    <RANKING order="3" place="3" resultid="2242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2237" />
                    <RANKING order="2" place="2" resultid="2242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="13" agemin="10" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2949" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1067" daytime="09:28" gender="M" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1068" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1663" />
                    <RANKING order="2" place="2" resultid="1444" />
                    <RANKING order="3" place="3" resultid="1658" />
                    <RANKING order="4" place="4" resultid="2252" />
                    <RANKING order="5" place="5" resultid="2256" />
                    <RANKING order="6" place="6" resultid="2246" />
                    <RANKING order="7" place="7" resultid="2688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1663" />
                    <RANKING order="2" place="2" resultid="1658" />
                    <RANKING order="3" place="3" resultid="2252" />
                    <RANKING order="4" place="4" resultid="2256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2246" />
                    <RANKING order="2" place="2" resultid="2688" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2950" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1071" daytime="09:34" gender="F" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1072" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1693" />
                    <RANKING order="2" place="2" resultid="2148" />
                    <RANKING order="3" place="3" resultid="2159" />
                    <RANKING order="4" place="4" resultid="2664" />
                    <RANKING order="5" place="5" resultid="2719" />
                    <RANKING order="6" place="6" resultid="1667" />
                    <RANKING order="7" place="7" resultid="1677" />
                    <RANKING order="8" place="8" resultid="1697" />
                    <RANKING order="9" place="9" resultid="1967" />
                    <RANKING order="10" place="10" resultid="2698" />
                    <RANKING order="11" place="11" resultid="1672" />
                    <RANKING order="12" place="11" resultid="2389" />
                    <RANKING order="13" place="13" resultid="2261" />
                    <RANKING order="14" place="14" resultid="2162" />
                    <RANKING order="15" place="15" resultid="1713" />
                    <RANKING order="16" place="16" resultid="2722" />
                    <RANKING order="17" place="17" resultid="1630" />
                    <RANKING order="18" place="18" resultid="2490" />
                    <RANKING order="19" place="19" resultid="1890" />
                    <RANKING order="20" place="20" resultid="2725" />
                    <RANKING order="21" place="21" resultid="1457" />
                    <RANKING order="22" place="22" resultid="2271" />
                    <RANKING order="23" place="23" resultid="2446" />
                    <RANKING order="24" place="24" resultid="2153" />
                    <RANKING order="25" place="24" resultid="2432" />
                    <RANKING order="26" place="26" resultid="1701" />
                    <RANKING order="27" place="27" resultid="2027" />
                    <RANKING order="28" place="28" resultid="2376" />
                    <RANKING order="29" place="29" resultid="1259" />
                    <RANKING order="30" place="30" resultid="1390" />
                    <RANKING order="31" place="31" resultid="2693" />
                    <RANKING order="32" place="32" resultid="1901" />
                    <RANKING order="33" place="33" resultid="2190" />
                    <RANKING order="34" place="34" resultid="2703" />
                    <RANKING order="35" place="35" resultid="1690" />
                    <RANKING order="36" place="36" resultid="2451" />
                    <RANKING order="37" place="37" resultid="2275" />
                    <RANKING order="38" place="38" resultid="1461" />
                    <RANKING order="39" place="39" resultid="1464" />
                    <RANKING order="40" place="40" resultid="2098" />
                    <RANKING order="41" place="41" resultid="2501" />
                    <RANKING order="42" place="42" resultid="2106" />
                    <RANKING order="43" place="43" resultid="1963" />
                    <RANKING order="44" place="44" resultid="1709" />
                    <RANKING order="45" place="45" resultid="1604" />
                    <RANKING order="46" place="46" resultid="1718" />
                    <RANKING order="47" place="47" resultid="2019" />
                    <RANKING order="48" place="48" resultid="1975" />
                    <RANKING order="49" place="49" resultid="1705" />
                    <RANKING order="50" place="50" resultid="2428" />
                    <RANKING order="51" place="51" resultid="1468" />
                    <RANKING order="52" place="52" resultid="1282" />
                    <RANKING order="53" place="53" resultid="1476" />
                    <RANKING order="54" place="54" resultid="1617" />
                    <RANKING order="55" place="55" resultid="1613" />
                    <RANKING order="56" place="56" resultid="2267" />
                    <RANKING order="57" place="57" resultid="2114" />
                    <RANKING order="58" place="58" resultid="1912" />
                    <RANKING order="59" place="59" resultid="1922" />
                    <RANKING order="60" place="60" resultid="2102" />
                    <RANKING order="61" place="61" resultid="2110" />
                    <RANKING order="62" place="62" resultid="1609" />
                    <RANKING order="63" place="63" resultid="1312" />
                    <RANKING order="64" place="64" resultid="1625" />
                    <RANKING order="65" place="65" resultid="1315" />
                    <RANKING order="66" place="66" resultid="1472" />
                    <RANKING order="67" place="67" resultid="1449" />
                    <RANKING order="68" place="68" resultid="1917" />
                    <RANKING order="69" place="69" resultid="1621" />
                    <RANKING order="70" place="70" resultid="1189" />
                    <RANKING order="71" place="71" resultid="2023" />
                    <RANKING order="72" place="72" resultid="2457" />
                    <RANKING order="73" place="73" resultid="1907" />
                    <RANKING order="74" place="74" resultid="1896" />
                    <RANKING order="75" place="75" resultid="1402" />
                    <RANKING order="76" place="76" resultid="3081" />
                    <RANKING order="77" place="77" resultid="2638" />
                    <RANKING order="78" place="78" resultid="1341" />
                    <RANKING order="79" place="79" resultid="2461" />
                    <RANKING order="80" place="80" resultid="1394" />
                    <RANKING order="81" place="81" resultid="1398" />
                    <RANKING order="82" place="82" resultid="2589" />
                    <RANKING order="83" place="83" resultid="2494" />
                    <RANKING order="84" place="84" resultid="1681" />
                    <RANKING order="85" place="85" resultid="2498" />
                    <RANKING order="86" place="86" resultid="1686" />
                    <RANKING order="87" place="-1" resultid="1212" />
                    <RANKING order="88" place="-1" resultid="1364" />
                    <RANKING order="89" place="-1" resultid="1452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2159" />
                    <RANKING order="2" place="2" resultid="2719" />
                    <RANKING order="3" place="3" resultid="1667" />
                    <RANKING order="4" place="4" resultid="1677" />
                    <RANKING order="5" place="5" resultid="2698" />
                    <RANKING order="6" place="6" resultid="1672" />
                    <RANKING order="7" place="6" resultid="2389" />
                    <RANKING order="8" place="8" resultid="2261" />
                    <RANKING order="9" place="9" resultid="1713" />
                    <RANKING order="10" place="10" resultid="2490" />
                    <RANKING order="11" place="11" resultid="1890" />
                    <RANKING order="12" place="12" resultid="2725" />
                    <RANKING order="13" place="13" resultid="2446" />
                    <RANKING order="14" place="14" resultid="2376" />
                    <RANKING order="15" place="15" resultid="1390" />
                    <RANKING order="16" place="16" resultid="2693" />
                    <RANKING order="17" place="17" resultid="1901" />
                    <RANKING order="18" place="18" resultid="2190" />
                    <RANKING order="19" place="19" resultid="2703" />
                    <RANKING order="20" place="20" resultid="1690" />
                    <RANKING order="21" place="21" resultid="2275" />
                    <RANKING order="22" place="22" resultid="1461" />
                    <RANKING order="23" place="23" resultid="1464" />
                    <RANKING order="24" place="24" resultid="1963" />
                    <RANKING order="25" place="25" resultid="1709" />
                    <RANKING order="26" place="26" resultid="1718" />
                    <RANKING order="27" place="27" resultid="2019" />
                    <RANKING order="28" place="28" resultid="1705" />
                    <RANKING order="29" place="29" resultid="1468" />
                    <RANKING order="30" place="30" resultid="1282" />
                    <RANKING order="31" place="31" resultid="1476" />
                    <RANKING order="32" place="32" resultid="1617" />
                    <RANKING order="33" place="33" resultid="2267" />
                    <RANKING order="34" place="34" resultid="1449" />
                    <RANKING order="35" place="35" resultid="1621" />
                    <RANKING order="36" place="36" resultid="1189" />
                    <RANKING order="37" place="37" resultid="1896" />
                    <RANKING order="38" place="38" resultid="1394" />
                    <RANKING order="39" place="-1" resultid="1364" />
                    <RANKING order="40" place="-1" resultid="1452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1967" />
                    <RANKING order="2" place="2" resultid="2451" />
                    <RANKING order="3" place="3" resultid="2098" />
                    <RANKING order="4" place="4" resultid="2106" />
                    <RANKING order="5" place="5" resultid="1604" />
                    <RANKING order="6" place="6" resultid="1975" />
                    <RANKING order="7" place="7" resultid="1613" />
                    <RANKING order="8" place="8" resultid="2114" />
                    <RANKING order="9" place="9" resultid="1912" />
                    <RANKING order="10" place="10" resultid="1922" />
                    <RANKING order="11" place="11" resultid="2102" />
                    <RANKING order="12" place="12" resultid="2110" />
                    <RANKING order="13" place="13" resultid="1609" />
                    <RANKING order="14" place="14" resultid="1625" />
                    <RANKING order="15" place="15" resultid="1472" />
                    <RANKING order="16" place="16" resultid="1917" />
                    <RANKING order="17" place="17" resultid="2023" />
                    <RANKING order="18" place="18" resultid="2457" />
                    <RANKING order="19" place="19" resultid="1907" />
                    <RANKING order="20" place="20" resultid="1402" />
                    <RANKING order="21" place="21" resultid="3081" />
                    <RANKING order="22" place="22" resultid="2638" />
                    <RANKING order="23" place="23" resultid="1341" />
                    <RANKING order="24" place="24" resultid="2461" />
                    <RANKING order="25" place="25" resultid="1398" />
                    <RANKING order="26" place="26" resultid="2589" />
                    <RANKING order="27" place="-1" resultid="1212" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2951" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2952" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2953" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2954" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2955" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2956" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2957" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="2958" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="2959" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" daytime="09:46" gender="M" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1076" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2806" />
                    <RANKING order="2" place="2" resultid="2669" />
                    <RANKING order="3" place="3" resultid="2728" />
                    <RANKING order="4" place="4" resultid="1726" />
                    <RANKING order="5" place="5" resultid="2732" />
                    <RANKING order="6" place="6" resultid="1294" />
                    <RANKING order="7" place="7" resultid="2290" />
                    <RANKING order="8" place="8" resultid="1415" />
                    <RANKING order="9" place="9" resultid="1331" />
                    <RANKING order="10" place="10" resultid="2004" />
                    <RANKING order="11" place="11" resultid="2745" />
                    <RANKING order="12" place="12" resultid="1488" />
                    <RANKING order="13" place="13" resultid="2597" />
                    <RANKING order="14" place="14" resultid="2592" />
                    <RANKING order="15" place="15" resultid="2065" />
                    <RANKING order="16" place="16" resultid="2436" />
                    <RANKING order="17" place="17" resultid="1327" />
                    <RANKING order="18" place="18" resultid="1721" />
                    <RANKING order="19" place="19" resultid="2674" />
                    <RANKING order="20" place="20" resultid="2060" />
                    <RANKING order="21" place="21" resultid="2740" />
                    <RANKING order="22" place="22" resultid="2736" />
                    <RANKING order="23" place="23" resultid="1506" />
                    <RANKING order="24" place="24" resultid="1749" />
                    <RANKING order="25" place="25" resultid="1765" />
                    <RANKING order="26" place="26" resultid="1929" />
                    <RANKING order="27" place="27" resultid="2226" />
                    <RANKING order="28" place="28" resultid="1637" />
                    <RANKING order="29" place="29" resultid="1984" />
                    <RANKING order="30" place="30" resultid="1276" />
                    <RANKING order="31" place="31" resultid="2605" />
                    <RANKING order="32" place="32" resultid="2510" />
                    <RANKING order="33" place="33" resultid="1290" />
                    <RANKING order="34" place="34" resultid="2708" />
                    <RANKING order="35" place="35" resultid="1510" />
                    <RANKING order="36" place="35" resultid="2613" />
                    <RANKING order="37" place="37" resultid="2609" />
                    <RANKING order="38" place="38" resultid="1493" />
                    <RANKING order="39" place="39" resultid="1501" />
                    <RANKING order="40" place="40" resultid="2030" />
                    <RANKING order="41" place="41" resultid="1514" />
                    <RANKING order="42" place="42" resultid="2601" />
                    <RANKING order="43" place="43" resultid="1286" />
                    <RANKING order="44" place="44" resultid="1760" />
                    <RANKING order="45" place="45" resultid="1754" />
                    <RANKING order="46" place="46" resultid="1498" />
                    <RANKING order="47" place="47" resultid="1771" />
                    <RANKING order="48" place="48" resultid="2514" />
                    <RANKING order="49" place="49" resultid="2194" />
                    <RANKING order="50" place="50" resultid="2118" />
                    <RANKING order="51" place="51" resultid="2531" />
                    <RANKING order="52" place="52" resultid="2535" />
                    <RANKING order="53" place="53" resultid="1528" />
                    <RANKING order="54" place="54" resultid="1979" />
                    <RANKING order="55" place="55" resultid="2523" />
                    <RANKING order="56" place="56" resultid="1484" />
                    <RANKING order="57" place="57" resultid="2200" />
                    <RANKING order="58" place="58" resultid="1191" />
                    <RANKING order="59" place="59" resultid="2465" />
                    <RANKING order="60" place="60" resultid="1757" />
                    <RANKING order="61" place="61" resultid="2143" />
                    <RANKING order="62" place="61" resultid="2469" />
                    <RANKING order="63" place="63" resultid="1406" />
                    <RANKING order="64" place="64" resultid="2049" />
                    <RANKING order="65" place="65" resultid="2505" />
                    <RANKING order="66" place="66" resultid="1523" />
                    <RANKING order="67" place="67" resultid="2285" />
                    <RANKING order="68" place="68" resultid="2041" />
                    <RANKING order="69" place="69" resultid="2038" />
                    <RANKING order="70" place="69" resultid="2415" />
                    <RANKING order="71" place="71" resultid="1989" />
                    <RANKING order="72" place="72" resultid="2473" />
                    <RANKING order="73" place="73" resultid="2407" />
                    <RANKING order="74" place="74" resultid="1481" />
                    <RANKING order="75" place="75" resultid="1642" />
                    <RANKING order="76" place="76" resultid="1538" />
                    <RANKING order="77" place="77" resultid="2945" />
                    <RANKING order="78" place="78" resultid="2518" />
                    <RANKING order="79" place="79" resultid="2395" />
                    <RANKING order="80" place="80" resultid="1647" />
                    <RANKING order="81" place="81" resultid="2034" />
                    <RANKING order="82" place="82" resultid="1734" />
                    <RANKING order="83" place="83" resultid="2477" />
                    <RANKING order="84" place="84" resultid="1739" />
                    <RANKING order="85" place="85" resultid="2527" />
                    <RANKING order="86" place="86" resultid="1217" />
                    <RANKING order="87" place="87" resultid="1195" />
                    <RANKING order="88" place="88" resultid="2618" />
                    <RANKING order="89" place="89" resultid="1934" />
                    <RANKING order="90" place="90" resultid="1633" />
                    <RANKING order="91" place="91" resultid="1411" />
                    <RANKING order="92" place="92" resultid="1744" />
                    <RANKING order="93" place="93" resultid="2481" />
                    <RANKING order="94" place="94" resultid="2045" />
                    <RANKING order="95" place="95" resultid="1319" />
                    <RANKING order="96" place="96" resultid="1940" />
                    <RANKING order="97" place="97" resultid="1996" />
                    <RANKING order="98" place="98" resultid="2053" />
                    <RANKING order="99" place="99" resultid="2365" />
                    <RANKING order="100" place="100" resultid="2000" />
                    <RANKING order="101" place="101" resultid="1193" />
                    <RANKING order="102" place="102" resultid="2280" />
                    <RANKING order="103" place="103" resultid="1344" />
                    <RANKING order="104" place="104" resultid="2008" />
                    <RANKING order="105" place="105" resultid="1222" />
                    <RANKING order="106" place="106" resultid="2139" />
                    <RANKING order="107" place="107" resultid="1729" />
                    <RANKING order="108" place="108" resultid="2412" />
                    <RANKING order="109" place="109" resultid="2643" />
                    <RANKING order="110" place="-1" resultid="1993" />
                    <RANKING order="111" place="-1" resultid="1368" />
                    <RANKING order="112" place="-1" resultid="1519" />
                    <RANKING order="113" place="-1" resultid="1533" />
                    <RANKING order="114" place="-1" resultid="1763" />
                    <RANKING order="115" place="-1" resultid="1769" />
                    <RANKING order="116" place="-1" resultid="2057" />
                    <RANKING order="117" place="-1" resultid="2123" />
                    <RANKING order="118" place="-1" resultid="2197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2669" />
                    <RANKING order="2" place="2" resultid="2745" />
                    <RANKING order="3" place="3" resultid="2065" />
                    <RANKING order="4" place="4" resultid="2436" />
                    <RANKING order="5" place="5" resultid="2674" />
                    <RANKING order="6" place="6" resultid="1765" />
                    <RANKING order="7" place="7" resultid="1929" />
                    <RANKING order="8" place="8" resultid="1637" />
                    <RANKING order="9" place="9" resultid="1984" />
                    <RANKING order="10" place="10" resultid="1276" />
                    <RANKING order="11" place="11" resultid="2605" />
                    <RANKING order="12" place="12" resultid="2708" />
                    <RANKING order="13" place="13" resultid="1510" />
                    <RANKING order="14" place="13" resultid="2613" />
                    <RANKING order="15" place="15" resultid="2030" />
                    <RANKING order="16" place="16" resultid="1514" />
                    <RANKING order="17" place="17" resultid="1286" />
                    <RANKING order="18" place="18" resultid="1760" />
                    <RANKING order="19" place="19" resultid="1498" />
                    <RANKING order="20" place="20" resultid="2514" />
                    <RANKING order="21" place="21" resultid="2194" />
                    <RANKING order="22" place="22" resultid="2531" />
                    <RANKING order="23" place="23" resultid="2535" />
                    <RANKING order="24" place="24" resultid="1528" />
                    <RANKING order="25" place="25" resultid="2523" />
                    <RANKING order="26" place="26" resultid="1484" />
                    <RANKING order="27" place="27" resultid="2200" />
                    <RANKING order="28" place="28" resultid="2465" />
                    <RANKING order="29" place="29" resultid="1757" />
                    <RANKING order="30" place="30" resultid="2469" />
                    <RANKING order="31" place="31" resultid="1406" />
                    <RANKING order="32" place="32" resultid="2049" />
                    <RANKING order="33" place="33" resultid="1523" />
                    <RANKING order="34" place="34" resultid="2041" />
                    <RANKING order="35" place="35" resultid="2038" />
                    <RANKING order="36" place="36" resultid="2473" />
                    <RANKING order="37" place="37" resultid="1481" />
                    <RANKING order="38" place="38" resultid="1642" />
                    <RANKING order="39" place="39" resultid="2518" />
                    <RANKING order="40" place="40" resultid="2034" />
                    <RANKING order="41" place="41" resultid="2477" />
                    <RANKING order="42" place="42" resultid="2527" />
                    <RANKING order="43" place="43" resultid="1195" />
                    <RANKING order="44" place="44" resultid="1633" />
                    <RANKING order="45" place="45" resultid="2481" />
                    <RANKING order="46" place="46" resultid="2045" />
                    <RANKING order="47" place="-1" resultid="1368" />
                    <RANKING order="48" place="-1" resultid="1519" />
                    <RANKING order="49" place="-1" resultid="2057" />
                    <RANKING order="50" place="-1" resultid="2197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1754" />
                    <RANKING order="2" place="2" resultid="2118" />
                    <RANKING order="3" place="3" resultid="1191" />
                    <RANKING order="4" place="4" resultid="2285" />
                    <RANKING order="5" place="5" resultid="1989" />
                    <RANKING order="6" place="6" resultid="1538" />
                    <RANKING order="7" place="7" resultid="2395" />
                    <RANKING order="8" place="8" resultid="1647" />
                    <RANKING order="9" place="9" resultid="1739" />
                    <RANKING order="10" place="10" resultid="1217" />
                    <RANKING order="11" place="11" resultid="2618" />
                    <RANKING order="12" place="12" resultid="1934" />
                    <RANKING order="13" place="13" resultid="1411" />
                    <RANKING order="14" place="14" resultid="1744" />
                    <RANKING order="15" place="15" resultid="1940" />
                    <RANKING order="16" place="16" resultid="1996" />
                    <RANKING order="17" place="17" resultid="2053" />
                    <RANKING order="18" place="18" resultid="2000" />
                    <RANKING order="19" place="19" resultid="1193" />
                    <RANKING order="20" place="20" resultid="2280" />
                    <RANKING order="21" place="21" resultid="1344" />
                    <RANKING order="22" place="22" resultid="2008" />
                    <RANKING order="23" place="23" resultid="1222" />
                    <RANKING order="24" place="24" resultid="2643" />
                    <RANKING order="25" place="-1" resultid="1993" />
                    <RANKING order="26" place="-1" resultid="1533" />
                    <RANKING order="27" place="-1" resultid="1763" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2960" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2961" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2962" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2963" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2964" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2965" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2966" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="2967" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="2968" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="2969" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="2970" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="2971" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1079" daytime="10:02" gender="F" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1420" />
                    <RANKING order="2" place="2" resultid="2748" />
                    <RANKING order="3" place="3" resultid="2379" />
                    <RANKING order="4" place="4" resultid="2069" />
                    <RANKING order="5" place="5" resultid="2028" />
                    <RANKING order="6" place="6" resultid="1307" />
                    <RANKING order="7" place="7" resultid="1423" />
                    <RANKING order="8" place="8" resultid="1777" />
                    <RANKING order="9" place="9" resultid="2652" />
                    <RANKING order="10" place="10" resultid="2485" />
                    <RANKING order="11" place="11" resultid="1431" />
                    <RANKING order="12" place="12" resultid="1226" />
                    <RANKING order="13" place="13" resultid="2621" />
                    <RANKING order="14" place="14" resultid="2011" />
                    <RANKING order="15" place="15" resultid="1427" />
                    <RANKING order="16" place="16" resultid="1682" />
                    <RANKING order="17" place="17" resultid="1775" />
                    <RANKING order="18" place="18" resultid="1687" />
                    <RANKING order="19" place="-1" resultid="1213" />
                    <RANKING order="20" place="-1" resultid="1543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1420" />
                    <RANKING order="2" place="2" resultid="2379" />
                    <RANKING order="3" place="3" resultid="2069" />
                    <RANKING order="4" place="4" resultid="1423" />
                    <RANKING order="5" place="-1" resultid="1543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1777" />
                    <RANKING order="2" place="2" resultid="2652" />
                    <RANKING order="3" place="3" resultid="2485" />
                    <RANKING order="4" place="4" resultid="1431" />
                    <RANKING order="5" place="5" resultid="1226" />
                    <RANKING order="6" place="6" resultid="2621" />
                    <RANKING order="7" place="7" resultid="2011" />
                    <RANKING order="8" place="8" resultid="1427" />
                    <RANKING order="9" place="-1" resultid="1213" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2972" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2973" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1083" daytime="10:12" gender="M" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1084" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1552" />
                    <RANKING order="2" place="2" resultid="1797" />
                    <RANKING order="3" place="3" resultid="2751" />
                    <RANKING order="4" place="4" resultid="2295" />
                    <RANKING order="5" place="5" resultid="2061" />
                    <RANKING order="6" place="6" resultid="1556" />
                    <RANKING order="7" place="7" resultid="1809" />
                    <RANKING order="8" place="8" resultid="1336" />
                    <RANKING order="9" place="9" resultid="1801" />
                    <RANKING order="10" place="10" resultid="1782" />
                    <RANKING order="11" place="11" resultid="1548" />
                    <RANKING order="12" place="12" resultid="2077" />
                    <RANKING order="13" place="13" resultid="2633" />
                    <RANKING order="14" place="14" resultid="2074" />
                    <RANKING order="15" place="15" resultid="1790" />
                    <RANKING order="16" place="16" resultid="2247" />
                    <RANKING order="17" place="17" resultid="2506" />
                    <RANKING order="18" place="18" resultid="1347" />
                    <RANKING order="19" place="19" resultid="2204" />
                    <RANKING order="20" place="20" resultid="1787" />
                    <RANKING order="21" place="21" resultid="2625" />
                    <RANKING order="22" place="22" resultid="1435" />
                    <RANKING order="23" place="23" resultid="2646" />
                    <RANKING order="24" place="24" resultid="1264" />
                    <RANKING order="25" place="25" resultid="1268" />
                    <RANKING order="26" place="-1" resultid="2257" />
                    <RANKING order="27" place="-1" resultid="2421" />
                    <RANKING order="28" place="-1" resultid="1793" />
                    <RANKING order="29" place="-1" resultid="1805" />
                    <RANKING order="30" place="-1" resultid="1351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2751" />
                    <RANKING order="2" place="2" resultid="1556" />
                    <RANKING order="3" place="3" resultid="1809" />
                    <RANKING order="4" place="4" resultid="1801" />
                    <RANKING order="5" place="5" resultid="1548" />
                    <RANKING order="6" place="6" resultid="2077" />
                    <RANKING order="7" place="7" resultid="2074" />
                    <RANKING order="8" place="8" resultid="1790" />
                    <RANKING order="9" place="-1" resultid="2257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2633" />
                    <RANKING order="2" place="2" resultid="2247" />
                    <RANKING order="3" place="3" resultid="1347" />
                    <RANKING order="4" place="4" resultid="2204" />
                    <RANKING order="5" place="5" resultid="2625" />
                    <RANKING order="6" place="6" resultid="1435" />
                    <RANKING order="7" place="7" resultid="2646" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2974" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2975" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2976" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1087" daytime="10:24" gender="F" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1088" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2665" />
                    <RANKING order="2" place="2" resultid="1816" />
                    <RANKING order="3" place="3" resultid="2761" />
                    <RANKING order="4" place="4" resultid="2758" />
                    <RANKING order="5" place="5" resultid="1668" />
                    <RANKING order="6" place="6" resultid="2679" />
                    <RANKING order="7" place="7" resultid="1260" />
                    <RANKING order="8" place="8" resultid="2262" />
                    <RANKING order="9" place="9" resultid="2154" />
                    <RANKING order="10" place="10" resultid="2163" />
                    <RANKING order="11" place="11" resultid="2302" />
                    <RANKING order="12" place="12" resultid="2390" />
                    <RANKING order="13" place="13" resultid="2082" />
                    <RANKING order="14" place="14" resultid="2764" />
                    <RANKING order="15" place="15" resultid="2755" />
                    <RANKING order="16" place="16" resultid="1453" />
                    <RANKING order="17" place="17" resultid="1813" />
                    <RANKING order="18" place="18" resultid="2694" />
                    <RANKING order="19" place="19" resultid="2452" />
                    <RANKING order="20" place="20" resultid="1567" />
                    <RANKING order="21" place="21" resultid="2298" />
                    <RANKING order="22" place="22" resultid="1560" />
                    <RANKING order="23" place="23" resultid="1563" />
                    <RANKING order="24" place="24" resultid="1945" />
                    <RANKING order="25" place="-1" resultid="1370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2761" />
                    <RANKING order="2" place="2" resultid="1668" />
                    <RANKING order="3" place="3" resultid="2262" />
                    <RANKING order="4" place="4" resultid="2302" />
                    <RANKING order="5" place="5" resultid="2390" />
                    <RANKING order="6" place="6" resultid="2082" />
                    <RANKING order="7" place="7" resultid="2764" />
                    <RANKING order="8" place="8" resultid="2755" />
                    <RANKING order="9" place="9" resultid="1453" />
                    <RANKING order="10" place="10" resultid="2694" />
                    <RANKING order="11" place="11" resultid="2298" />
                    <RANKING order="12" place="12" resultid="1560" />
                    <RANKING order="13" place="-1" resultid="1370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1813" />
                    <RANKING order="2" place="2" resultid="2452" />
                    <RANKING order="3" place="3" resultid="1567" />
                    <RANKING order="4" place="4" resultid="1563" />
                    <RANKING order="5" place="5" resultid="1945" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2977" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2978" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2979" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1091" daytime="10:30" gender="M" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1092" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1823" />
                    <RANKING order="2" place="2" resultid="1416" />
                    <RANKING order="3" place="3" resultid="1576" />
                    <RANKING order="4" place="4" resultid="2768" />
                    <RANKING order="5" place="5" resultid="2670" />
                    <RANKING order="6" place="6" resultid="2310" />
                    <RANKING order="7" place="7" resultid="2675" />
                    <RANKING order="8" place="8" resultid="2086" />
                    <RANKING order="9" place="9" resultid="1291" />
                    <RANKING order="10" place="10" resultid="1255" />
                    <RANKING order="11" place="11" resultid="1502" />
                    <RANKING order="12" place="12" resultid="1298" />
                    <RANKING order="13" place="13" resultid="2539" />
                    <RANKING order="14" place="14" resultid="1277" />
                    <RANKING order="15" place="15" resultid="2306" />
                    <RANKING order="16" place="16" resultid="2709" />
                    <RANKING order="17" place="17" resultid="1197" />
                    <RANKING order="18" place="18" resultid="2089" />
                    <RANKING order="19" place="19" resultid="1571" />
                    <RANKING order="20" place="20" resultid="2078" />
                    <RANKING order="21" place="21" resultid="2416" />
                    <RANKING order="22" place="22" resultid="2810" />
                    <RANKING order="23" place="23" resultid="1580" />
                    <RANKING order="24" place="24" resultid="1412" />
                    <RANKING order="25" place="25" resultid="1539" />
                    <RANKING order="26" place="26" resultid="1820" />
                    <RANKING order="27" place="27" resultid="2127" />
                    <RANKING order="28" place="28" resultid="2629" />
                    <RANKING order="29" place="29" resultid="2713" />
                    <RANKING order="30" place="30" resultid="1382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2670" />
                    <RANKING order="2" place="2" resultid="2675" />
                    <RANKING order="3" place="3" resultid="2086" />
                    <RANKING order="4" place="4" resultid="1298" />
                    <RANKING order="5" place="5" resultid="2539" />
                    <RANKING order="6" place="6" resultid="1277" />
                    <RANKING order="7" place="7" resultid="2306" />
                    <RANKING order="8" place="8" resultid="2709" />
                    <RANKING order="9" place="9" resultid="1197" />
                    <RANKING order="10" place="10" resultid="2089" />
                    <RANKING order="11" place="11" resultid="2078" />
                    <RANKING order="12" place="12" resultid="2810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1580" />
                    <RANKING order="2" place="2" resultid="1412" />
                    <RANKING order="3" place="3" resultid="1539" />
                    <RANKING order="4" place="4" resultid="2629" />
                    <RANKING order="5" place="5" resultid="2713" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2980" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2981" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2982" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1095" daytime="10:38" gender="F" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1096" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2683" />
                    <RANKING order="2" place="2" resultid="2149" />
                    <RANKING order="3" place="3" resultid="1826" />
                    <RANKING order="4" place="4" resultid="1714" />
                    <RANKING order="5" place="5" resultid="2765" />
                    <RANKING order="6" place="6" resultid="2371" />
                    <RANKING order="7" place="7" resultid="1673" />
                    <RANKING order="8" place="8" resultid="1828" />
                    <RANKING order="9" place="9" resultid="2319" />
                    <RANKING order="10" place="10" resultid="2447" />
                    <RANKING order="11" place="11" resultid="2391" />
                    <RANKING order="12" place="12" resultid="2327" />
                    <RANKING order="13" place="13" resultid="2243" />
                    <RANKING order="14" place="14" resultid="2323" />
                    <RANKING order="15" place="15" resultid="2212" />
                    <RANKING order="16" place="16" resultid="2433" />
                    <RANKING order="17" place="17" resultid="2233" />
                    <RANKING order="18" place="18" resultid="2502" />
                    <RANKING order="19" place="19" resultid="2704" />
                    <RANKING order="20" place="20" resultid="2299" />
                    <RANKING order="21" place="21" resultid="2331" />
                    <RANKING order="22" place="22" resultid="2020" />
                    <RANKING order="23" place="23" resultid="1477" />
                    <RANKING order="24" place="24" resultid="1918" />
                    <RANKING order="25" place="25" resultid="1949" />
                    <RANKING order="26" place="26" resultid="1923" />
                    <RANKING order="27" place="27" resultid="2314" />
                    <RANKING order="28" place="28" resultid="2115" />
                    <RANKING order="29" place="29" resultid="2103" />
                    <RANKING order="30" place="30" resultid="1622" />
                    <RANKING order="31" place="31" resultid="1954" />
                    <RANKING order="32" place="32" resultid="2024" />
                    <RANKING order="33" place="33" resultid="1913" />
                    <RANKING order="34" place="34" resultid="1908" />
                    <RANKING order="35" place="35" resultid="1395" />
                    <RANKING order="36" place="36" resultid="2462" />
                    <RANKING order="37" place="37" resultid="1399" />
                    <RANKING order="38" place="38" resultid="2543" />
                    <RANKING order="39" place="-1" resultid="1891" />
                    <RANKING order="40" place="-1" resultid="1365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1826" />
                    <RANKING order="2" place="2" resultid="1714" />
                    <RANKING order="3" place="3" resultid="2765" />
                    <RANKING order="4" place="4" resultid="2371" />
                    <RANKING order="5" place="5" resultid="1673" />
                    <RANKING order="6" place="6" resultid="2447" />
                    <RANKING order="7" place="7" resultid="2391" />
                    <RANKING order="8" place="8" resultid="2327" />
                    <RANKING order="9" place="9" resultid="2243" />
                    <RANKING order="10" place="10" resultid="2323" />
                    <RANKING order="11" place="11" resultid="2212" />
                    <RANKING order="12" place="12" resultid="2704" />
                    <RANKING order="13" place="13" resultid="2299" />
                    <RANKING order="14" place="14" resultid="2331" />
                    <RANKING order="15" place="15" resultid="2020" />
                    <RANKING order="16" place="16" resultid="1477" />
                    <RANKING order="17" place="17" resultid="2314" />
                    <RANKING order="18" place="18" resultid="1622" />
                    <RANKING order="19" place="19" resultid="1395" />
                    <RANKING order="20" place="-1" resultid="1891" />
                    <RANKING order="21" place="-1" resultid="1365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1918" />
                    <RANKING order="2" place="2" resultid="1949" />
                    <RANKING order="3" place="3" resultid="1923" />
                    <RANKING order="4" place="4" resultid="2115" />
                    <RANKING order="5" place="5" resultid="2103" />
                    <RANKING order="6" place="6" resultid="1954" />
                    <RANKING order="7" place="7" resultid="2024" />
                    <RANKING order="8" place="8" resultid="1913" />
                    <RANKING order="9" place="9" resultid="1908" />
                    <RANKING order="10" place="10" resultid="2462" />
                    <RANKING order="11" place="11" resultid="1399" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2983" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2984" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2985" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2986" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2987" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1099" daytime="10:48" gender="M" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1100" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2733" />
                    <RANKING order="2" place="2" resultid="2774" />
                    <RANKING order="3" place="3" resultid="2729" />
                    <RANKING order="4" place="4" resultid="2593" />
                    <RANKING order="5" place="5" resultid="1838" />
                    <RANKING order="6" place="6" resultid="2778" />
                    <RANKING order="7" place="7" resultid="1507" />
                    <RANKING order="8" place="8" resultid="1295" />
                    <RANKING order="9" place="9" resultid="2005" />
                    <RANKING order="10" place="10" resultid="2781" />
                    <RANKING order="11" place="11" resultid="2253" />
                    <RANKING order="12" place="12" resultid="2741" />
                    <RANKING order="13" place="13" resultid="1236" />
                    <RANKING order="14" place="14" resultid="1659" />
                    <RANKING order="15" place="15" resultid="1766" />
                    <RANKING order="16" place="16" resultid="1849" />
                    <RANKING order="17" place="17" resultid="2291" />
                    <RANKING order="18" place="18" resultid="2550" />
                    <RANKING order="19" place="19" resultid="1332" />
                    <RANKING order="20" place="20" resultid="1515" />
                    <RANKING order="21" place="21" resultid="2227" />
                    <RANKING order="22" place="22" resultid="1930" />
                    <RANKING order="23" place="23" resultid="1489" />
                    <RANKING order="24" place="24" resultid="2657" />
                    <RANKING order="25" place="25" resultid="2540" />
                    <RANKING order="26" place="26" resultid="1833" />
                    <RANKING order="27" place="27" resultid="2532" />
                    <RANKING order="28" place="28" resultid="1842" />
                    <RANKING order="29" place="29" resultid="1524" />
                    <RANKING order="30" place="30" resultid="2385" />
                    <RANKING order="31" place="31" resultid="1355" />
                    <RANKING order="32" place="32" resultid="1846" />
                    <RANKING order="33" place="33" resultid="2470" />
                    <RANKING order="34" place="34" resultid="1643" />
                    <RANKING order="35" place="35" resultid="1585" />
                    <RANKING order="36" place="36" resultid="2286" />
                    <RANKING order="37" place="37" resultid="2216" />
                    <RANKING order="38" place="37" resultid="2408" />
                    <RANKING order="39" place="39" resultid="2546" />
                    <RANKING order="40" place="40" resultid="2050" />
                    <RANKING order="41" place="41" resultid="1200" />
                    <RANKING order="42" place="42" resultid="1581" />
                    <RANKING order="43" place="43" resultid="2396" />
                    <RANKING order="44" place="44" resultid="1997" />
                    <RANKING order="45" place="45" resultid="2689" />
                    <RANKING order="46" place="46" resultid="1218" />
                    <RANKING order="47" place="47" resultid="2046" />
                    <RANKING order="48" place="48" resultid="1634" />
                    <RANKING order="49" place="49" resultid="1345" />
                    <RANKING order="50" place="50" resultid="2366" />
                    <RANKING order="51" place="51" resultid="2554" />
                    <RANKING order="52" place="52" resultid="2561" />
                    <RANKING order="53" place="53" resultid="1223" />
                    <RANKING order="54" place="54" resultid="2281" />
                    <RANKING order="55" place="55" resultid="1730" />
                    <RANKING order="56" place="56" resultid="2558" />
                    <RANKING order="57" place="-1" resultid="1375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1838" />
                    <RANKING order="2" place="2" resultid="2253" />
                    <RANKING order="3" place="3" resultid="1236" />
                    <RANKING order="4" place="4" resultid="1659" />
                    <RANKING order="5" place="5" resultid="1766" />
                    <RANKING order="6" place="6" resultid="2550" />
                    <RANKING order="7" place="7" resultid="1515" />
                    <RANKING order="8" place="8" resultid="1930" />
                    <RANKING order="9" place="9" resultid="2657" />
                    <RANKING order="10" place="10" resultid="2540" />
                    <RANKING order="11" place="11" resultid="2532" />
                    <RANKING order="12" place="12" resultid="1842" />
                    <RANKING order="13" place="13" resultid="1524" />
                    <RANKING order="14" place="14" resultid="2385" />
                    <RANKING order="15" place="15" resultid="1846" />
                    <RANKING order="16" place="16" resultid="2470" />
                    <RANKING order="17" place="17" resultid="1643" />
                    <RANKING order="18" place="18" resultid="1585" />
                    <RANKING order="19" place="19" resultid="2546" />
                    <RANKING order="20" place="20" resultid="2050" />
                    <RANKING order="21" place="21" resultid="2046" />
                    <RANKING order="22" place="22" resultid="1634" />
                    <RANKING order="23" place="-1" resultid="1375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2286" />
                    <RANKING order="2" place="2" resultid="2216" />
                    <RANKING order="3" place="3" resultid="1200" />
                    <RANKING order="4" place="4" resultid="1581" />
                    <RANKING order="5" place="5" resultid="2396" />
                    <RANKING order="6" place="6" resultid="1997" />
                    <RANKING order="7" place="7" resultid="2689" />
                    <RANKING order="8" place="8" resultid="1218" />
                    <RANKING order="9" place="9" resultid="1345" />
                    <RANKING order="10" place="10" resultid="1223" />
                    <RANKING order="11" place="11" resultid="2281" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2988" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2989" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2990" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2991" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2992" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2993" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" daytime="10:58" gender="F" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1104" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1858" />
                    <RANKING order="2" place="2" resultid="2759" />
                    <RANKING order="3" place="3" resultid="2723" />
                    <RANKING order="4" place="4" resultid="2785" />
                    <RANKING order="5" place="5" resultid="2788" />
                    <RANKING order="6" place="6" resultid="1698" />
                    <RANKING order="7" place="7" resultid="2726" />
                    <RANKING order="8" place="8" resultid="2155" />
                    <RANKING order="9" place="9" resultid="1829" />
                    <RANKING order="10" place="10" resultid="1439" />
                    <RANKING order="11" place="11" resultid="2167" />
                    <RANKING order="12" place="12" resultid="1968" />
                    <RANKING order="13" place="13" resultid="2338" />
                    <RANKING order="14" place="14" resultid="1702" />
                    <RANKING order="15" place="15" resultid="2328" />
                    <RANKING order="16" place="16" resultid="2272" />
                    <RANKING order="17" place="17" resultid="2335" />
                    <RANKING order="18" place="18" resultid="2564" />
                    <RANKING order="19" place="19" resultid="1710" />
                    <RANKING order="20" place="20" resultid="1469" />
                    <RANKING order="21" place="21" resultid="1706" />
                    <RANKING order="22" place="22" resultid="2131" />
                    <RANKING order="23" place="23" resultid="1360" />
                    <RANKING order="24" place="24" resultid="1605" />
                    <RANKING order="25" place="25" resultid="2653" />
                    <RANKING order="26" place="26" resultid="1240" />
                    <RANKING order="27" place="27" resultid="2315" />
                    <RANKING order="28" place="28" resultid="1316" />
                    <RANKING order="29" place="29" resultid="1561" />
                    <RANKING order="30" place="30" resultid="1357" />
                    <RANKING order="31" place="31" resultid="1853" />
                    <RANKING order="32" place="-1" resultid="1371" />
                    <RANKING order="33" place="-1" resultid="1964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2785" />
                    <RANKING order="2" place="2" resultid="2726" />
                    <RANKING order="3" place="3" resultid="1439" />
                    <RANKING order="4" place="4" resultid="2167" />
                    <RANKING order="5" place="5" resultid="2338" />
                    <RANKING order="6" place="6" resultid="2328" />
                    <RANKING order="7" place="7" resultid="1710" />
                    <RANKING order="8" place="8" resultid="1469" />
                    <RANKING order="9" place="9" resultid="1706" />
                    <RANKING order="10" place="10" resultid="2315" />
                    <RANKING order="11" place="11" resultid="1561" />
                    <RANKING order="12" place="-1" resultid="1371" />
                    <RANKING order="13" place="-1" resultid="1964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1968" />
                    <RANKING order="2" place="2" resultid="2564" />
                    <RANKING order="3" place="3" resultid="1360" />
                    <RANKING order="4" place="4" resultid="1605" />
                    <RANKING order="5" place="5" resultid="2653" />
                    <RANKING order="6" place="6" resultid="1240" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2994" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2995" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2996" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2997" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="11:12" gender="M" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1445" />
                    <RANKING order="2" place="2" resultid="2343" />
                    <RANKING order="3" place="3" resultid="1866" />
                    <RANKING order="4" place="4" resultid="2511" />
                    <RANKING order="5" place="5" resultid="1590" />
                    <RANKING order="6" place="6" resultid="1244" />
                    <RANKING order="7" place="7" resultid="1494" />
                    <RANKING order="8" place="7" resultid="1870" />
                    <RANKING order="9" place="9" resultid="1572" />
                    <RANKING order="10" place="10" resultid="1772" />
                    <RANKING order="11" place="11" resultid="1985" />
                    <RANKING order="12" place="12" resultid="1722" />
                    <RANKING order="13" place="13" resultid="2572" />
                    <RANKING order="14" place="14" resultid="1549" />
                    <RANKING order="15" place="15" resultid="2606" />
                    <RANKING order="16" place="16" resultid="2031" />
                    <RANKING order="17" place="17" resultid="2536" />
                    <RANKING order="18" place="18" resultid="1980" />
                    <RANKING order="19" place="19" resultid="2602" />
                    <RANKING order="20" place="20" resultid="1511" />
                    <RANKING order="21" place="21" resultid="1407" />
                    <RANKING order="22" place="22" resultid="2575" />
                    <RANKING order="23" place="23" resultid="1862" />
                    <RANKING order="24" place="24" resultid="1529" />
                    <RANKING order="25" place="25" resultid="2248" />
                    <RANKING order="26" place="26" resultid="2035" />
                    <RANKING order="27" place="27" resultid="1219" />
                    <RANKING order="28" place="28" resultid="1735" />
                    <RANKING order="29" place="29" resultid="2690" />
                    <RANKING order="30" place="30" resultid="1247" />
                    <RANKING order="31" place="31" resultid="2578" />
                    <RANKING order="32" place="32" resultid="1821" />
                    <RANKING order="33" place="33" resultid="1383" />
                    <RANKING order="34" place="34" resultid="1323" />
                    <RANKING order="35" place="35" resultid="1303" />
                    <RANKING order="36" place="-1" resultid="1376" />
                    <RANKING order="37" place="-1" resultid="2124" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1590" />
                    <RANKING order="2" place="2" resultid="1244" />
                    <RANKING order="3" place="3" resultid="1985" />
                    <RANKING order="4" place="4" resultid="1549" />
                    <RANKING order="5" place="5" resultid="2606" />
                    <RANKING order="6" place="6" resultid="2031" />
                    <RANKING order="7" place="7" resultid="2536" />
                    <RANKING order="8" place="8" resultid="1511" />
                    <RANKING order="9" place="9" resultid="1407" />
                    <RANKING order="10" place="10" resultid="2575" />
                    <RANKING order="11" place="11" resultid="1529" />
                    <RANKING order="12" place="12" resultid="2035" />
                    <RANKING order="13" place="-1" resultid="1376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2248" />
                    <RANKING order="2" place="2" resultid="1219" />
                    <RANKING order="3" place="3" resultid="2690" />
                    <RANKING order="4" place="4" resultid="1247" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2998" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2999" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3000" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3001" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1111" daytime="11:26" gender="F" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1112" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2791" />
                    <RANKING order="2" place="2" resultid="1421" />
                    <RANKING order="3" place="3" resultid="2320" />
                    <RANKING order="4" place="4" resultid="2380" />
                    <RANKING order="5" place="5" resultid="2680" />
                    <RANKING order="6" place="6" resultid="1308" />
                    <RANKING order="7" place="7" resultid="2699" />
                    <RANKING order="8" place="8" resultid="1465" />
                    <RANKING order="9" place="9" resultid="1458" />
                    <RANKING order="10" place="10" resultid="2070" />
                    <RANKING order="11" place="11" resultid="1874" />
                    <RANKING order="12" place="12" resultid="1424" />
                    <RANKING order="13" place="13" resultid="1902" />
                    <RANKING order="14" place="14" resultid="1594" />
                    <RANKING order="15" place="15" resultid="1778" />
                    <RANKING order="16" place="16" resultid="2429" />
                    <RANKING order="17" place="17" resultid="2486" />
                    <RANKING order="18" place="18" resultid="2012" />
                    <RANKING order="19" place="19" resultid="1432" />
                    <RANKING order="20" place="20" resultid="1897" />
                    <RANKING order="21" place="21" resultid="2622" />
                    <RANKING order="22" place="22" resultid="1203" />
                    <RANKING order="23" place="23" resultid="1914" />
                    <RANKING order="24" place="24" resultid="1227" />
                    <RANKING order="25" place="25" resultid="1428" />
                    <RANKING order="26" place="26" resultid="2639" />
                    <RANKING order="27" place="27" resultid="1403" />
                    <RANKING order="28" place="28" resultid="1683" />
                    <RANKING order="29" place="29" resultid="1688" />
                    <RANKING order="30" place="-1" resultid="1214" />
                    <RANKING order="31" place="-1" resultid="1544" />
                    <RANKING order="32" place="-1" resultid="2268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2791" />
                    <RANKING order="2" place="2" resultid="1421" />
                    <RANKING order="3" place="3" resultid="2380" />
                    <RANKING order="4" place="4" resultid="2699" />
                    <RANKING order="5" place="5" resultid="1465" />
                    <RANKING order="6" place="6" resultid="2070" />
                    <RANKING order="7" place="7" resultid="1424" />
                    <RANKING order="8" place="8" resultid="1902" />
                    <RANKING order="9" place="9" resultid="1594" />
                    <RANKING order="10" place="10" resultid="1897" />
                    <RANKING order="11" place="-1" resultid="1544" />
                    <RANKING order="12" place="-1" resultid="2268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1874" />
                    <RANKING order="2" place="2" resultid="1778" />
                    <RANKING order="3" place="3" resultid="2486" />
                    <RANKING order="4" place="4" resultid="2012" />
                    <RANKING order="5" place="5" resultid="1432" />
                    <RANKING order="6" place="6" resultid="2622" />
                    <RANKING order="7" place="7" resultid="1203" />
                    <RANKING order="8" place="8" resultid="1914" />
                    <RANKING order="9" place="9" resultid="1227" />
                    <RANKING order="10" place="10" resultid="1428" />
                    <RANKING order="11" place="11" resultid="2639" />
                    <RANKING order="12" place="12" resultid="1403" />
                    <RANKING order="13" place="-1" resultid="1214" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3002" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3003" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3004" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3005" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1115" daytime="11:36" gender="M" number="15" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1116" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2598" />
                    <RANKING order="2" place="2" resultid="1750" />
                    <RANKING order="3" place="3" resultid="2797" />
                    <RANKING order="4" place="4" resultid="1553" />
                    <RANKING order="5" place="5" resultid="2794" />
                    <RANKING order="6" place="6" resultid="2782" />
                    <RANKING order="7" place="7" resultid="2258" />
                    <RANKING order="8" place="8" resultid="2066" />
                    <RANKING order="9" place="9" resultid="2752" />
                    <RANKING order="10" place="10" resultid="2170" />
                    <RANKING order="11" place="11" resultid="1557" />
                    <RANKING order="12" place="12" resultid="1798" />
                    <RANKING order="13" place="13" resultid="1877" />
                    <RANKING order="14" place="14" resultid="2062" />
                    <RANKING order="15" place="15" resultid="1783" />
                    <RANKING order="16" place="16" resultid="1802" />
                    <RANKING order="17" place="17" resultid="2676" />
                    <RANKING order="18" place="18" resultid="1810" />
                    <RANKING order="19" place="19" resultid="1337" />
                    <RANKING order="20" place="20" resultid="2800" />
                    <RANKING order="21" place="21" resultid="2092" />
                    <RANKING order="22" place="22" resultid="2075" />
                    <RANKING order="23" place="23" resultid="1299" />
                    <RANKING order="24" place="24" resultid="2079" />
                    <RANKING order="25" place="25" resultid="2634" />
                    <RANKING order="26" place="26" resultid="2610" />
                    <RANKING order="27" place="27" resultid="2042" />
                    <RANKING order="28" place="28" resultid="2507" />
                    <RANKING order="29" place="29" resultid="2582" />
                    <RANKING order="30" place="30" resultid="2519" />
                    <RANKING order="31" place="31" resultid="1352" />
                    <RANKING order="32" place="32" resultid="1348" />
                    <RANKING order="33" place="33" resultid="2482" />
                    <RANKING order="34" place="34" resultid="1788" />
                    <RANKING order="35" place="35" resultid="2422" />
                    <RANKING order="36" place="36" resultid="1941" />
                    <RANKING order="37" place="37" resultid="1740" />
                    <RANKING order="38" place="38" resultid="1206" />
                    <RANKING order="39" place="39" resultid="1436" />
                    <RANKING order="40" place="40" resultid="1248" />
                    <RANKING order="41" place="41" resultid="1320" />
                    <RANKING order="42" place="42" resultid="2647" />
                    <RANKING order="43" place="43" resultid="1265" />
                    <RANKING order="44" place="44" resultid="1935" />
                    <RANKING order="45" place="45" resultid="2714" />
                    <RANKING order="46" place="46" resultid="1269" />
                    <RANKING order="47" place="-1" resultid="1520" />
                    <RANKING order="48" place="-1" resultid="1534" />
                    <RANKING order="49" place="-1" resultid="1794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2258" />
                    <RANKING order="2" place="2" resultid="2066" />
                    <RANKING order="3" place="3" resultid="2752" />
                    <RANKING order="4" place="4" resultid="2170" />
                    <RANKING order="5" place="5" resultid="1557" />
                    <RANKING order="6" place="6" resultid="1877" />
                    <RANKING order="7" place="7" resultid="1802" />
                    <RANKING order="8" place="8" resultid="2676" />
                    <RANKING order="9" place="9" resultid="1810" />
                    <RANKING order="10" place="10" resultid="2800" />
                    <RANKING order="11" place="11" resultid="2092" />
                    <RANKING order="12" place="12" resultid="2075" />
                    <RANKING order="13" place="13" resultid="1299" />
                    <RANKING order="14" place="14" resultid="2079" />
                    <RANKING order="15" place="15" resultid="2042" />
                    <RANKING order="16" place="16" resultid="2519" />
                    <RANKING order="17" place="17" resultid="2482" />
                    <RANKING order="18" place="-1" resultid="1520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2634" />
                    <RANKING order="2" place="2" resultid="1348" />
                    <RANKING order="3" place="3" resultid="1941" />
                    <RANKING order="4" place="4" resultid="1740" />
                    <RANKING order="5" place="5" resultid="1206" />
                    <RANKING order="6" place="6" resultid="1436" />
                    <RANKING order="7" place="7" resultid="1248" />
                    <RANKING order="8" place="8" resultid="2647" />
                    <RANKING order="9" place="9" resultid="1935" />
                    <RANKING order="10" place="10" resultid="2714" />
                    <RANKING order="11" place="-1" resultid="1534" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3006" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3007" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3008" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3009" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3010" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1119" daytime="11:46" gender="F" number="16" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1120" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1694" />
                    <RANKING order="2" place="2" resultid="2666" />
                    <RANKING order="3" place="3" resultid="2150" />
                    <RANKING order="4" place="4" resultid="2238" />
                    <RANKING order="5" place="5" resultid="1669" />
                    <RANKING order="6" place="6" resultid="2766" />
                    <RANKING order="7" place="7" resultid="1678" />
                    <RANKING order="8" place="8" resultid="1674" />
                    <RANKING order="9" place="9" resultid="1892" />
                    <RANKING order="10" place="10" resultid="1817" />
                    <RANKING order="11" place="11" resultid="2762" />
                    <RANKING order="12" place="12" resultid="2263" />
                    <RANKING order="13" place="13" resultid="2392" />
                    <RANKING order="14" place="14" resultid="1261" />
                    <RANKING order="15" place="15" resultid="2303" />
                    <RANKING order="16" place="16" resultid="2209" />
                    <RANKING order="17" place="17" resultid="2156" />
                    <RANKING order="18" place="17" resultid="2448" />
                    <RANKING order="19" place="19" resultid="2244" />
                    <RANKING order="20" place="20" resultid="2491" />
                    <RANKING order="21" place="21" resultid="2352" />
                    <RANKING order="22" place="22" resultid="2276" />
                    <RANKING order="23" place="23" resultid="1454" />
                    <RANKING order="24" place="24" resultid="2695" />
                    <RANKING order="25" place="25" resultid="2213" />
                    <RANKING order="26" place="26" resultid="1814" />
                    <RANKING order="27" place="27" resultid="2565" />
                    <RANKING order="28" place="28" resultid="2453" />
                    <RANKING order="29" place="29" resultid="1568" />
                    <RANKING order="30" place="30" resultid="2332" />
                    <RANKING order="31" place="31" resultid="2339" />
                    <RANKING order="32" place="32" resultid="2107" />
                    <RANKING order="33" place="33" resultid="1903" />
                    <RANKING order="34" place="34" resultid="2300" />
                    <RANKING order="35" place="35" resultid="1976" />
                    <RANKING order="36" place="36" resultid="1283" />
                    <RANKING order="37" place="37" resultid="1924" />
                    <RANKING order="38" place="38" resultid="1618" />
                    <RANKING order="39" place="39" resultid="1919" />
                    <RANKING order="40" place="40" resultid="1950" />
                    <RANKING order="41" place="41" resultid="1626" />
                    <RANKING order="42" place="42" resultid="2441" />
                    <RANKING order="43" place="43" resultid="1473" />
                    <RANKING order="44" place="44" resultid="1946" />
                    <RANKING order="45" place="45" resultid="1955" />
                    <RANKING order="46" place="46" resultid="1564" />
                    <RANKING order="47" place="47" resultid="1909" />
                    <RANKING order="48" place="48" resultid="1342" />
                    <RANKING order="49" place="49" resultid="2463" />
                    <RANKING order="50" place="50" resultid="2495" />
                    <RANKING order="51" place="51" resultid="2499" />
                    <RANKING order="52" place="-1" resultid="1372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2238" />
                    <RANKING order="2" place="2" resultid="1669" />
                    <RANKING order="3" place="3" resultid="2766" />
                    <RANKING order="4" place="4" resultid="1678" />
                    <RANKING order="5" place="5" resultid="1674" />
                    <RANKING order="6" place="6" resultid="1892" />
                    <RANKING order="7" place="7" resultid="2762" />
                    <RANKING order="8" place="8" resultid="2263" />
                    <RANKING order="9" place="9" resultid="2392" />
                    <RANKING order="10" place="10" resultid="2303" />
                    <RANKING order="11" place="11" resultid="2209" />
                    <RANKING order="12" place="12" resultid="2448" />
                    <RANKING order="13" place="13" resultid="2244" />
                    <RANKING order="14" place="14" resultid="2491" />
                    <RANKING order="15" place="15" resultid="2352" />
                    <RANKING order="16" place="16" resultid="2276" />
                    <RANKING order="17" place="17" resultid="1454" />
                    <RANKING order="18" place="18" resultid="2695" />
                    <RANKING order="19" place="19" resultid="2213" />
                    <RANKING order="20" place="20" resultid="2332" />
                    <RANKING order="21" place="21" resultid="2339" />
                    <RANKING order="22" place="22" resultid="1903" />
                    <RANKING order="23" place="23" resultid="2300" />
                    <RANKING order="24" place="24" resultid="1283" />
                    <RANKING order="25" place="25" resultid="1618" />
                    <RANKING order="26" place="26" resultid="2441" />
                    <RANKING order="27" place="-1" resultid="1372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1814" />
                    <RANKING order="2" place="2" resultid="2565" />
                    <RANKING order="3" place="3" resultid="2453" />
                    <RANKING order="4" place="4" resultid="1568" />
                    <RANKING order="5" place="5" resultid="2107" />
                    <RANKING order="6" place="6" resultid="1976" />
                    <RANKING order="7" place="7" resultid="1924" />
                    <RANKING order="8" place="8" resultid="1919" />
                    <RANKING order="9" place="9" resultid="1950" />
                    <RANKING order="10" place="10" resultid="1626" />
                    <RANKING order="11" place="11" resultid="1473" />
                    <RANKING order="12" place="12" resultid="1946" />
                    <RANKING order="13" place="13" resultid="1955" />
                    <RANKING order="14" place="14" resultid="1564" />
                    <RANKING order="15" place="15" resultid="1909" />
                    <RANKING order="16" place="16" resultid="1342" />
                    <RANKING order="17" place="17" resultid="2463" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3011" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3012" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3013" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3014" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3015" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3016" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1123" daytime="11:56" gender="M" number="17" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1124" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1824" />
                    <RANKING order="2" place="2" resultid="2734" />
                    <RANKING order="3" place="3" resultid="2807" />
                    <RANKING order="4" place="4" resultid="2775" />
                    <RANKING order="5" place="5" resultid="2671" />
                    <RANKING order="6" place="6" resultid="2798" />
                    <RANKING order="7" place="7" resultid="1333" />
                    <RANKING order="8" place="8" resultid="2006" />
                    <RANKING order="9" place="9" resultid="1839" />
                    <RANKING order="10" place="10" resultid="1328" />
                    <RANKING order="11" place="11" resultid="1577" />
                    <RANKING order="12" place="12" resultid="1417" />
                    <RANKING order="13" place="13" resultid="2173" />
                    <RANKING order="14" place="14" resultid="2292" />
                    <RANKING order="15" place="15" resultid="2087" />
                    <RANKING order="16" place="16" resultid="2737" />
                    <RANKING order="17" place="17" resultid="2311" />
                    <RANKING order="18" place="18" resultid="2437" />
                    <RANKING order="19" place="19" resultid="1503" />
                    <RANKING order="20" place="20" resultid="1723" />
                    <RANKING order="21" place="21" resultid="1490" />
                    <RANKING order="22" place="22" resultid="1292" />
                    <RANKING order="23" place="23" resultid="2176" />
                    <RANKING order="24" place="24" resultid="2614" />
                    <RANKING order="25" place="25" resultid="2603" />
                    <RANKING order="26" place="26" resultid="1638" />
                    <RANKING order="27" place="27" resultid="2710" />
                    <RANKING order="28" place="28" resultid="2228" />
                    <RANKING order="29" place="29" resultid="2307" />
                    <RANKING order="30" place="30" resultid="1931" />
                    <RANKING order="31" place="31" resultid="1573" />
                    <RANKING order="32" place="32" resultid="1198" />
                    <RANKING order="33" place="33" resultid="1881" />
                    <RANKING order="34" place="34" resultid="2195" />
                    <RANKING order="35" place="35" resultid="2611" />
                    <RANKING order="36" place="36" resultid="2417" />
                    <RANKING order="37" place="37" resultid="2541" />
                    <RANKING order="38" place="38" resultid="1525" />
                    <RANKING order="39" place="39" resultid="2144" />
                    <RANKING order="40" place="40" resultid="2533" />
                    <RANKING order="41" place="41" resultid="1843" />
                    <RANKING order="42" place="42" resultid="1990" />
                    <RANKING order="43" place="43" resultid="2515" />
                    <RANKING order="44" place="43" resultid="2524" />
                    <RANKING order="45" place="45" resultid="1485" />
                    <RANKING order="46" place="46" resultid="1287" />
                    <RANKING order="47" place="47" resultid="2222" />
                    <RANKING order="48" place="48" resultid="2287" />
                    <RANKING order="49" place="49" resultid="2466" />
                    <RANKING order="50" place="50" resultid="2201" />
                    <RANKING order="51" place="51" resultid="2205" />
                    <RANKING order="52" place="52" resultid="1530" />
                    <RANKING order="53" place="53" resultid="1272" />
                    <RANKING order="54" place="54" resultid="1540" />
                    <RANKING order="55" place="55" resultid="1644" />
                    <RANKING order="56" place="56" resultid="2471" />
                    <RANKING order="57" place="57" resultid="1648" />
                    <RANKING order="58" place="57" resultid="1736" />
                    <RANKING order="59" place="59" resultid="2409" />
                    <RANKING order="60" place="60" resultid="2630" />
                    <RANKING order="61" place="61" resultid="2219" />
                    <RANKING order="62" place="62" resultid="2397" />
                    <RANKING order="63" place="63" resultid="2478" />
                    <RANKING order="64" place="64" resultid="2128" />
                    <RANKING order="65" place="65" resultid="2474" />
                    <RANKING order="66" place="66" resultid="2198" />
                    <RANKING order="67" place="67" resultid="2015" />
                    <RANKING order="68" place="68" resultid="2001" />
                    <RANKING order="69" place="69" resultid="1936" />
                    <RANKING order="70" place="70" resultid="2715" />
                    <RANKING order="71" place="71" resultid="2367" />
                    <RANKING order="72" place="72" resultid="2282" />
                    <RANKING order="73" place="73" resultid="2559" />
                    <RANKING order="74" place="-1" resultid="1582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2671" />
                    <RANKING order="2" place="2" resultid="1839" />
                    <RANKING order="3" place="3" resultid="2173" />
                    <RANKING order="4" place="4" resultid="2087" />
                    <RANKING order="5" place="5" resultid="2437" />
                    <RANKING order="6" place="6" resultid="2614" />
                    <RANKING order="7" place="7" resultid="1638" />
                    <RANKING order="8" place="8" resultid="2710" />
                    <RANKING order="9" place="9" resultid="2307" />
                    <RANKING order="10" place="10" resultid="1931" />
                    <RANKING order="11" place="11" resultid="1198" />
                    <RANKING order="12" place="12" resultid="1881" />
                    <RANKING order="13" place="13" resultid="2195" />
                    <RANKING order="14" place="14" resultid="2541" />
                    <RANKING order="15" place="15" resultid="1525" />
                    <RANKING order="16" place="16" resultid="2533" />
                    <RANKING order="17" place="17" resultid="1843" />
                    <RANKING order="18" place="18" resultid="2515" />
                    <RANKING order="19" place="18" resultid="2524" />
                    <RANKING order="20" place="20" resultid="1485" />
                    <RANKING order="21" place="21" resultid="1287" />
                    <RANKING order="22" place="22" resultid="2466" />
                    <RANKING order="23" place="23" resultid="2201" />
                    <RANKING order="24" place="24" resultid="1530" />
                    <RANKING order="25" place="25" resultid="1644" />
                    <RANKING order="26" place="26" resultid="2471" />
                    <RANKING order="27" place="27" resultid="2219" />
                    <RANKING order="28" place="28" resultid="2478" />
                    <RANKING order="29" place="29" resultid="2474" />
                    <RANKING order="30" place="30" resultid="2198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1990" />
                    <RANKING order="2" place="2" resultid="2222" />
                    <RANKING order="3" place="3" resultid="2287" />
                    <RANKING order="4" place="4" resultid="2205" />
                    <RANKING order="5" place="5" resultid="1540" />
                    <RANKING order="6" place="6" resultid="1648" />
                    <RANKING order="7" place="7" resultid="2630" />
                    <RANKING order="8" place="8" resultid="2397" />
                    <RANKING order="9" place="9" resultid="2015" />
                    <RANKING order="10" place="10" resultid="2001" />
                    <RANKING order="11" place="11" resultid="1936" />
                    <RANKING order="12" place="12" resultid="2715" />
                    <RANKING order="13" place="13" resultid="2282" />
                    <RANKING order="14" place="-1" resultid="1582" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3017" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3018" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3019" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3020" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3021" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3022" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="3023" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="3024" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1127" daytime="13:00" gender="F" number="18" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1128" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1715" />
                    <RANKING order="2" place="2" resultid="2372" />
                    <RANKING order="3" place="3" resultid="1830" />
                    <RANKING order="4" place="4" resultid="2324" />
                    <RANKING order="5" place="5" resultid="1597" />
                    <RANKING order="6" place="6" resultid="2705" />
                    <RANKING order="7" place="7" resultid="2099" />
                    <RANKING order="8" place="8" resultid="1241" />
                    <RANKING order="9" place="9" resultid="2316" />
                    <RANKING order="10" place="10" resultid="3082" />
                    <RANKING order="11" place="11" resultid="1478" />
                    <RANKING order="12" place="12" resultid="1854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1715" />
                    <RANKING order="2" place="2" resultid="2372" />
                    <RANKING order="3" place="3" resultid="2324" />
                    <RANKING order="4" place="4" resultid="1597" />
                    <RANKING order="5" place="5" resultid="2705" />
                    <RANKING order="6" place="6" resultid="2316" />
                    <RANKING order="7" place="7" resultid="1478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2099" />
                    <RANKING order="2" place="2" resultid="1241" />
                    <RANKING order="3" place="3" resultid="3082" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3025" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3026" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1131" daytime="13:08" gender="M" number="19" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1132" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1278" />
                    <RANKING order="2" place="2" resultid="1591" />
                    <RANKING order="3" place="3" resultid="1237" />
                    <RANKING order="4" place="4" resultid="2386" />
                    <RANKING order="5" place="5" resultid="2249" />
                    <RANKING order="6" place="6" resultid="1586" />
                    <RANKING order="7" place="7" resultid="1834" />
                    <RANKING order="8" place="8" resultid="2217" />
                    <RANKING order="9" place="9" resultid="2223" />
                    <RANKING order="10" place="10" resultid="2691" />
                    <RANKING order="11" place="11" resultid="2423" />
                    <RANKING order="12" place="12" resultid="2585" />
                    <RANKING order="13" place="13" resultid="2555" />
                    <RANKING order="14" place="-1" resultid="1377" />
                    <RANKING order="15" place="-1" resultid="1850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1133" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1278" />
                    <RANKING order="2" place="2" resultid="1591" />
                    <RANKING order="3" place="3" resultid="1237" />
                    <RANKING order="4" place="4" resultid="2386" />
                    <RANKING order="5" place="5" resultid="1586" />
                    <RANKING order="6" place="-1" resultid="1377" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2249" />
                    <RANKING order="2" place="2" resultid="2217" />
                    <RANKING order="3" place="3" resultid="2223" />
                    <RANKING order="4" place="4" resultid="2691" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3027" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3028" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" daytime="13:16" gender="F" number="20" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1136" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1695" />
                    <RANKING order="2" place="2" resultid="1859" />
                    <RANKING order="3" place="3" resultid="2160" />
                    <RANKING order="4" place="4" resultid="2749" />
                    <RANKING order="5" place="5" resultid="2720" />
                    <RANKING order="6" place="6" resultid="1670" />
                    <RANKING order="7" place="7" resultid="1631" />
                    <RANKING order="8" place="8" resultid="1699" />
                    <RANKING order="9" place="9" resultid="2264" />
                    <RANKING order="10" place="10" resultid="2234" />
                    <RANKING order="11" place="11" resultid="2179" />
                    <RANKING order="12" place="12" resultid="2164" />
                    <RANKING order="13" place="13" resultid="2700" />
                    <RANKING order="14" place="14" resultid="2393" />
                    <RANKING order="15" place="15" resultid="2157" />
                    <RANKING order="16" place="16" resultid="2329" />
                    <RANKING order="17" place="17" resultid="1440" />
                    <RANKING order="18" place="18" resultid="1893" />
                    <RANKING order="19" place="19" resultid="1703" />
                    <RANKING order="20" place="20" resultid="2277" />
                    <RANKING order="21" place="21" resultid="1391" />
                    <RANKING order="22" place="22" resultid="2340" />
                    <RANKING order="23" place="23" resultid="2191" />
                    <RANKING order="24" place="24" resultid="1904" />
                    <RANKING order="25" place="25" resultid="1691" />
                    <RANKING order="26" place="26" resultid="2503" />
                    <RANKING order="27" place="27" resultid="1711" />
                    <RANKING order="28" place="28" resultid="1462" />
                    <RANKING order="29" place="29" resultid="2108" />
                    <RANKING order="30" place="29" resultid="2696" />
                    <RANKING order="31" place="31" resultid="2100" />
                    <RANKING order="32" place="32" resultid="1707" />
                    <RANKING order="33" place="33" resultid="1719" />
                    <RANKING order="34" place="34" resultid="1606" />
                    <RANKING order="35" place="35" resultid="2654" />
                    <RANKING order="36" place="36" resultid="2269" />
                    <RANKING order="37" place="37" resultid="1569" />
                    <RANKING order="38" place="38" resultid="1614" />
                    <RANKING order="39" place="39" resultid="1313" />
                    <RANKING order="40" place="40" resultid="1619" />
                    <RANKING order="41" place="41" resultid="2111" />
                    <RANKING order="42" place="42" resultid="1610" />
                    <RANKING order="43" place="43" resultid="1474" />
                    <RANKING order="44" place="44" resultid="1317" />
                    <RANKING order="45" place="45" resultid="2116" />
                    <RANKING order="46" place="46" resultid="1925" />
                    <RANKING order="47" place="47" resultid="1627" />
                    <RANKING order="48" place="48" resultid="2104" />
                    <RANKING order="49" place="49" resultid="2025" />
                    <RANKING order="50" place="50" resultid="2458" />
                    <RANKING order="51" place="51" resultid="1898" />
                    <RANKING order="52" place="52" resultid="1450" />
                    <RANKING order="53" place="53" resultid="1956" />
                    <RANKING order="54" place="54" resultid="1947" />
                    <RANKING order="55" place="55" resultid="1565" />
                    <RANKING order="56" place="56" resultid="1855" />
                    <RANKING order="57" place="57" resultid="2640" />
                    <RANKING order="58" place="-1" resultid="1366" />
                    <RANKING order="59" place="-1" resultid="1373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2160" />
                    <RANKING order="2" place="2" resultid="2720" />
                    <RANKING order="3" place="3" resultid="1670" />
                    <RANKING order="4" place="4" resultid="2264" />
                    <RANKING order="5" place="5" resultid="2700" />
                    <RANKING order="6" place="6" resultid="2393" />
                    <RANKING order="7" place="7" resultid="2329" />
                    <RANKING order="8" place="8" resultid="1440" />
                    <RANKING order="9" place="9" resultid="1893" />
                    <RANKING order="10" place="10" resultid="2277" />
                    <RANKING order="11" place="11" resultid="1391" />
                    <RANKING order="12" place="12" resultid="2340" />
                    <RANKING order="13" place="13" resultid="2191" />
                    <RANKING order="14" place="14" resultid="1904" />
                    <RANKING order="15" place="15" resultid="1691" />
                    <RANKING order="16" place="16" resultid="1711" />
                    <RANKING order="17" place="17" resultid="1462" />
                    <RANKING order="18" place="18" resultid="2696" />
                    <RANKING order="19" place="19" resultid="1707" />
                    <RANKING order="20" place="20" resultid="1719" />
                    <RANKING order="21" place="21" resultid="2269" />
                    <RANKING order="22" place="22" resultid="1619" />
                    <RANKING order="23" place="23" resultid="1898" />
                    <RANKING order="24" place="24" resultid="1450" />
                    <RANKING order="25" place="-1" resultid="1366" />
                    <RANKING order="26" place="-1" resultid="1373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2108" />
                    <RANKING order="2" place="2" resultid="2100" />
                    <RANKING order="3" place="3" resultid="1606" />
                    <RANKING order="4" place="4" resultid="2654" />
                    <RANKING order="5" place="5" resultid="1569" />
                    <RANKING order="6" place="6" resultid="1614" />
                    <RANKING order="7" place="7" resultid="2111" />
                    <RANKING order="8" place="8" resultid="1610" />
                    <RANKING order="9" place="9" resultid="1474" />
                    <RANKING order="10" place="10" resultid="2116" />
                    <RANKING order="11" place="11" resultid="1925" />
                    <RANKING order="12" place="12" resultid="1627" />
                    <RANKING order="13" place="13" resultid="2104" />
                    <RANKING order="14" place="14" resultid="2025" />
                    <RANKING order="15" place="15" resultid="2458" />
                    <RANKING order="16" place="16" resultid="1956" />
                    <RANKING order="17" place="17" resultid="1947" />
                    <RANKING order="18" place="18" resultid="1565" />
                    <RANKING order="19" place="19" resultid="2640" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3029" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3030" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3031" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3032" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3033" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3034" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1139" daytime="13:28" gender="M" number="21" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1140" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1418" />
                    <RANKING order="2" place="1" resultid="2808" />
                    <RANKING order="3" place="3" resultid="2594" />
                    <RANKING order="4" place="4" resultid="2672" />
                    <RANKING order="5" place="5" resultid="2344" />
                    <RANKING order="6" place="6" resultid="2067" />
                    <RANKING order="7" place="7" resultid="2803" />
                    <RANKING order="8" place="8" resultid="1446" />
                    <RANKING order="9" place="9" resultid="1840" />
                    <RANKING order="10" place="10" resultid="1867" />
                    <RANKING order="11" place="11" resultid="2746" />
                    <RANKING order="12" place="12" resultid="1724" />
                    <RANKING order="13" place="13" resultid="2182" />
                    <RANKING order="14" place="14" resultid="1329" />
                    <RANKING order="15" place="15" resultid="2742" />
                    <RANKING order="16" place="16" resultid="1491" />
                    <RANKING order="17" place="17" resultid="2438" />
                    <RANKING order="18" place="18" resultid="2512" />
                    <RANKING order="19" place="19" resultid="2174" />
                    <RANKING order="20" place="20" resultid="1574" />
                    <RANKING order="21" place="21" resultid="2738" />
                    <RANKING order="22" place="22" resultid="1495" />
                    <RANKING order="23" place="23" resultid="1932" />
                    <RANKING order="24" place="24" resultid="2177" />
                    <RANKING order="25" place="25" resultid="1871" />
                    <RANKING order="26" place="26" resultid="1592" />
                    <RANKING order="27" place="27" resultid="2615" />
                    <RANKING order="28" place="28" resultid="2711" />
                    <RANKING order="29" place="29" resultid="2607" />
                    <RANKING order="30" place="30" resultid="1550" />
                    <RANKING order="31" place="31" resultid="2032" />
                    <RANKING order="32" place="32" resultid="1773" />
                    <RANKING order="33" place="33" resultid="1639" />
                    <RANKING order="34" place="34" resultid="2516" />
                    <RANKING order="35" place="35" resultid="1755" />
                    <RANKING order="36" place="36" resultid="1512" />
                    <RANKING order="37" place="37" resultid="1882" />
                    <RANKING order="38" place="38" resultid="2658" />
                    <RANKING order="39" place="39" resultid="2525" />
                    <RANKING order="40" place="40" resultid="1758" />
                    <RANKING order="41" place="41" resultid="2119" />
                    <RANKING order="42" place="42" resultid="1981" />
                    <RANKING order="43" place="43" resultid="2467" />
                    <RANKING order="44" place="44" resultid="1499" />
                    <RANKING order="45" place="45" resultid="1408" />
                    <RANKING order="46" place="46" resultid="2145" />
                    <RANKING order="47" place="47" resultid="2039" />
                    <RANKING order="48" place="48" resultid="2418" />
                    <RANKING order="49" place="49" resultid="2090" />
                    <RANKING order="50" place="50" resultid="2051" />
                    <RANKING order="51" place="51" resultid="2520" />
                    <RANKING order="52" place="52" resultid="2508" />
                    <RANKING order="53" place="53" resultid="1531" />
                    <RANKING order="54" place="54" resultid="2547" />
                    <RANKING order="55" place="55" resultid="1482" />
                    <RANKING order="56" place="56" resultid="1541" />
                    <RANKING order="57" place="57" resultid="2528" />
                    <RANKING order="58" place="58" resultid="2579" />
                    <RANKING order="59" place="59" resultid="2036" />
                    <RANKING order="60" place="60" resultid="2220" />
                    <RANKING order="61" place="61" resultid="1220" />
                    <RANKING order="62" place="62" resultid="2479" />
                    <RANKING order="63" place="63" resultid="1413" />
                    <RANKING order="64" place="64" resultid="1937" />
                    <RANKING order="65" place="65" resultid="1635" />
                    <RANKING order="66" place="66" resultid="2047" />
                    <RANKING order="67" place="67" resultid="1994" />
                    <RANKING order="68" place="68" resultid="2619" />
                    <RANKING order="69" place="69" resultid="1745" />
                    <RANKING order="70" place="70" resultid="1942" />
                    <RANKING order="71" place="71" resultid="2054" />
                    <RANKING order="72" place="72" resultid="2016" />
                    <RANKING order="73" place="73" resultid="2002" />
                    <RANKING order="74" place="74" resultid="2368" />
                    <RANKING order="75" place="75" resultid="2009" />
                    <RANKING order="76" place="76" resultid="1731" />
                    <RANKING order="77" place="-1" resultid="1288" />
                    <RANKING order="78" place="-1" resultid="1296" />
                    <RANKING order="79" place="-1" resultid="1535" />
                    <RANKING order="80" place="-1" resultid="1806" />
                    <RANKING order="81" place="-1" resultid="2058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1141" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2672" />
                    <RANKING order="2" place="2" resultid="2067" />
                    <RANKING order="3" place="3" resultid="2803" />
                    <RANKING order="4" place="4" resultid="1840" />
                    <RANKING order="5" place="5" resultid="2746" />
                    <RANKING order="6" place="6" resultid="2182" />
                    <RANKING order="7" place="7" resultid="2438" />
                    <RANKING order="8" place="8" resultid="2174" />
                    <RANKING order="9" place="9" resultid="1932" />
                    <RANKING order="10" place="10" resultid="1592" />
                    <RANKING order="11" place="11" resultid="2615" />
                    <RANKING order="12" place="12" resultid="2711" />
                    <RANKING order="13" place="13" resultid="2607" />
                    <RANKING order="14" place="14" resultid="1550" />
                    <RANKING order="15" place="15" resultid="2032" />
                    <RANKING order="16" place="16" resultid="1639" />
                    <RANKING order="17" place="17" resultid="2516" />
                    <RANKING order="18" place="18" resultid="1512" />
                    <RANKING order="19" place="19" resultid="1882" />
                    <RANKING order="20" place="20" resultid="2658" />
                    <RANKING order="21" place="21" resultid="2525" />
                    <RANKING order="22" place="22" resultid="1758" />
                    <RANKING order="23" place="23" resultid="2467" />
                    <RANKING order="24" place="24" resultid="1499" />
                    <RANKING order="25" place="25" resultid="1408" />
                    <RANKING order="26" place="26" resultid="2039" />
                    <RANKING order="27" place="27" resultid="2090" />
                    <RANKING order="28" place="28" resultid="2051" />
                    <RANKING order="29" place="29" resultid="2520" />
                    <RANKING order="30" place="30" resultid="1531" />
                    <RANKING order="31" place="31" resultid="2547" />
                    <RANKING order="32" place="32" resultid="1482" />
                    <RANKING order="33" place="33" resultid="2528" />
                    <RANKING order="34" place="34" resultid="2036" />
                    <RANKING order="35" place="35" resultid="2220" />
                    <RANKING order="36" place="36" resultid="2479" />
                    <RANKING order="37" place="37" resultid="1635" />
                    <RANKING order="38" place="38" resultid="2047" />
                    <RANKING order="39" place="-1" resultid="1288" />
                    <RANKING order="40" place="-1" resultid="2058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1755" />
                    <RANKING order="2" place="2" resultid="2119" />
                    <RANKING order="3" place="3" resultid="1541" />
                    <RANKING order="4" place="4" resultid="1220" />
                    <RANKING order="5" place="5" resultid="1413" />
                    <RANKING order="6" place="6" resultid="1937" />
                    <RANKING order="7" place="7" resultid="1994" />
                    <RANKING order="8" place="8" resultid="2619" />
                    <RANKING order="9" place="9" resultid="1745" />
                    <RANKING order="10" place="10" resultid="1942" />
                    <RANKING order="11" place="11" resultid="2054" />
                    <RANKING order="12" place="12" resultid="2016" />
                    <RANKING order="13" place="13" resultid="2002" />
                    <RANKING order="14" place="14" resultid="2009" />
                    <RANKING order="15" place="-1" resultid="1535" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3035" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3036" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3037" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3038" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3039" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3040" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="3041" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="3042" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="3043" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1143" daytime="13:46" gender="F" number="22" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1144" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2321" />
                    <RANKING order="2" place="2" resultid="2701" />
                    <RANKING order="3" place="3" resultid="2239" />
                    <RANKING order="4" place="4" resultid="2151" />
                    <RANKING order="5" place="5" resultid="1459" />
                    <RANKING order="6" place="6" resultid="2681" />
                    <RANKING order="7" place="7" resultid="2786" />
                    <RANKING order="8" place="8" resultid="2353" />
                    <RANKING order="9" place="9" resultid="1675" />
                    <RANKING order="10" place="10" resultid="1309" />
                    <RANKING order="11" place="11" resultid="2210" />
                    <RANKING order="12" place="12" resultid="1466" />
                    <RANKING order="13" place="13" resultid="2071" />
                    <RANKING order="14" place="14" resultid="2492" />
                    <RANKING order="15" place="15" resultid="1969" />
                    <RANKING order="16" place="16" resultid="1875" />
                    <RANKING order="17" place="17" resultid="2273" />
                    <RANKING order="18" place="18" resultid="1425" />
                    <RANKING order="19" place="19" resultid="1905" />
                    <RANKING order="20" place="20" resultid="1595" />
                    <RANKING order="21" place="21" resultid="1779" />
                    <RANKING order="22" place="22" resultid="2655" />
                    <RANKING order="23" place="23" resultid="2021" />
                    <RANKING order="24" place="24" resultid="2487" />
                    <RANKING order="25" place="25" resultid="2430" />
                    <RANKING order="26" place="26" resultid="2566" />
                    <RANKING order="27" place="27" resultid="2454" />
                    <RANKING order="28" place="28" resultid="1470" />
                    <RANKING order="29" place="29" resultid="2317" />
                    <RANKING order="30" place="30" resultid="1915" />
                    <RANKING order="31" place="31" resultid="2013" />
                    <RANKING order="32" place="32" resultid="1433" />
                    <RANKING order="33" place="33" resultid="1204" />
                    <RANKING order="34" place="34" resultid="1951" />
                    <RANKING order="35" place="35" resultid="2442" />
                    <RANKING order="36" place="36" resultid="2459" />
                    <RANKING order="37" place="37" resultid="1899" />
                    <RANKING order="38" place="38" resultid="2112" />
                    <RANKING order="39" place="39" resultid="1228" />
                    <RANKING order="40" place="40" resultid="1429" />
                    <RANKING order="41" place="41" resultid="1926" />
                    <RANKING order="42" place="42" resultid="1396" />
                    <RANKING order="43" place="43" resultid="1920" />
                    <RANKING order="44" place="44" resultid="2641" />
                    <RANKING order="45" place="45" resultid="1404" />
                    <RANKING order="46" place="46" resultid="1400" />
                    <RANKING order="47" place="47" resultid="1684" />
                    <RANKING order="48" place="48" resultid="2590" />
                    <RANKING order="49" place="49" resultid="2544" />
                    <RANKING order="50" place="-1" resultid="1215" />
                    <RANKING order="51" place="-1" resultid="1284" />
                    <RANKING order="52" place="-1" resultid="1545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2701" />
                    <RANKING order="2" place="2" resultid="2239" />
                    <RANKING order="3" place="3" resultid="2786" />
                    <RANKING order="4" place="4" resultid="2353" />
                    <RANKING order="5" place="5" resultid="1675" />
                    <RANKING order="6" place="6" resultid="2210" />
                    <RANKING order="7" place="7" resultid="1466" />
                    <RANKING order="8" place="8" resultid="2071" />
                    <RANKING order="9" place="9" resultid="2492" />
                    <RANKING order="10" place="10" resultid="1425" />
                    <RANKING order="11" place="11" resultid="1905" />
                    <RANKING order="12" place="12" resultid="1595" />
                    <RANKING order="13" place="13" resultid="2021" />
                    <RANKING order="14" place="14" resultid="1470" />
                    <RANKING order="15" place="15" resultid="2317" />
                    <RANKING order="16" place="16" resultid="2442" />
                    <RANKING order="17" place="17" resultid="1899" />
                    <RANKING order="18" place="18" resultid="1396" />
                    <RANKING order="19" place="-1" resultid="1284" />
                    <RANKING order="20" place="-1" resultid="1545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1969" />
                    <RANKING order="2" place="2" resultid="1875" />
                    <RANKING order="3" place="3" resultid="1779" />
                    <RANKING order="4" place="4" resultid="2655" />
                    <RANKING order="5" place="5" resultid="2487" />
                    <RANKING order="6" place="6" resultid="2566" />
                    <RANKING order="7" place="7" resultid="2454" />
                    <RANKING order="8" place="8" resultid="1915" />
                    <RANKING order="9" place="9" resultid="2013" />
                    <RANKING order="10" place="10" resultid="1433" />
                    <RANKING order="11" place="11" resultid="1204" />
                    <RANKING order="12" place="12" resultid="1951" />
                    <RANKING order="13" place="13" resultid="2459" />
                    <RANKING order="14" place="14" resultid="2112" />
                    <RANKING order="15" place="15" resultid="1228" />
                    <RANKING order="16" place="16" resultid="1429" />
                    <RANKING order="17" place="17" resultid="1926" />
                    <RANKING order="18" place="18" resultid="1920" />
                    <RANKING order="19" place="19" resultid="2641" />
                    <RANKING order="20" place="20" resultid="1404" />
                    <RANKING order="21" place="21" resultid="1400" />
                    <RANKING order="22" place="22" resultid="2590" />
                    <RANKING order="23" place="-1" resultid="1215" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3044" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3045" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3046" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3047" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3048" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3049" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1147" daytime="13:56" gender="M" number="23" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1148" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2599" />
                    <RANKING order="2" place="2" resultid="1554" />
                    <RANKING order="3" place="3" resultid="2783" />
                    <RANKING order="4" place="4" resultid="1751" />
                    <RANKING order="5" place="5" resultid="2753" />
                    <RANKING order="6" place="6" resultid="1664" />
                    <RANKING order="7" place="7" resultid="1558" />
                    <RANKING order="8" place="8" resultid="2171" />
                    <RANKING order="9" place="9" resultid="1799" />
                    <RANKING order="10" place="10" resultid="2801" />
                    <RANKING order="11" place="11" resultid="1784" />
                    <RANKING order="12" place="12" resultid="1334" />
                    <RANKING order="13" place="13" resultid="2063" />
                    <RANKING order="14" place="14" resultid="1660" />
                    <RANKING order="15" place="15" resultid="2229" />
                    <RANKING order="16" place="16" resultid="1803" />
                    <RANKING order="17" place="17" resultid="1878" />
                    <RANKING order="18" place="18" resultid="1761" />
                    <RANKING order="19" place="19" resultid="2293" />
                    <RANKING order="20" place="20" resultid="1986" />
                    <RANKING order="21" place="21" resultid="2677" />
                    <RANKING order="22" place="22" resultid="2776" />
                    <RANKING order="23" place="23" resultid="2093" />
                    <RANKING order="24" place="24" resultid="1811" />
                    <RANKING order="25" place="25" resultid="2551" />
                    <RANKING order="26" place="26" resultid="1516" />
                    <RANKING order="27" place="27" resultid="2080" />
                    <RANKING order="28" place="28" resultid="2548" />
                    <RANKING order="29" place="29" resultid="1486" />
                    <RANKING order="30" place="30" resultid="1844" />
                    <RANKING order="31" place="31" resultid="2635" />
                    <RANKING order="32" place="32" resultid="2659" />
                    <RANKING order="33" place="33" resultid="2043" />
                    <RANKING order="34" place="34" resultid="1791" />
                    <RANKING order="35" place="35" resultid="2583" />
                    <RANKING order="36" place="36" resultid="1349" />
                    <RANKING order="37" place="37" resultid="2202" />
                    <RANKING order="38" place="38" resultid="1353" />
                    <RANKING order="39" place="39" resultid="2521" />
                    <RANKING order="40" place="40" resultid="1209" />
                    <RANKING order="41" place="41" resultid="2288" />
                    <RANKING order="42" place="42" resultid="2626" />
                    <RANKING order="43" place="43" resultid="2475" />
                    <RANKING order="44" place="44" resultid="2483" />
                    <RANKING order="45" place="45" resultid="2129" />
                    <RANKING order="46" place="46" resultid="1587" />
                    <RANKING order="47" place="47" resultid="1649" />
                    <RANKING order="48" place="48" resultid="1943" />
                    <RANKING order="49" place="49" resultid="1437" />
                    <RANKING order="50" place="50" resultid="1741" />
                    <RANKING order="51" place="51" resultid="1266" />
                    <RANKING order="52" place="52" resultid="1207" />
                    <RANKING order="53" place="53" resultid="2134" />
                    <RANKING order="54" place="54" resultid="1938" />
                    <RANKING order="55" place="55" resultid="2529" />
                    <RANKING order="56" place="56" resultid="1321" />
                    <RANKING order="57" place="57" resultid="2398" />
                    <RANKING order="58" place="58" resultid="2136" />
                    <RANKING order="59" place="59" resultid="1249" />
                    <RANKING order="60" place="60" resultid="1746" />
                    <RANKING order="61" place="61" resultid="2648" />
                    <RANKING order="62" place="62" resultid="2716" />
                    <RANKING order="63" place="63" resultid="2055" />
                    <RANKING order="64" place="64" resultid="2140" />
                    <RANKING order="65" place="65" resultid="1224" />
                    <RANKING order="66" place="66" resultid="1270" />
                    <RANKING order="67" place="67" resultid="2644" />
                    <RANKING order="68" place="-1" resultid="1300" />
                    <RANKING order="69" place="-1" resultid="1521" />
                    <RANKING order="70" place="-1" resultid="1536" />
                    <RANKING order="71" place="-1" resultid="1795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1149" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2753" />
                    <RANKING order="2" place="2" resultid="1664" />
                    <RANKING order="3" place="3" resultid="1558" />
                    <RANKING order="4" place="4" resultid="2171" />
                    <RANKING order="5" place="5" resultid="2801" />
                    <RANKING order="6" place="6" resultid="1660" />
                    <RANKING order="7" place="7" resultid="1803" />
                    <RANKING order="8" place="8" resultid="1878" />
                    <RANKING order="9" place="9" resultid="1761" />
                    <RANKING order="10" place="10" resultid="1986" />
                    <RANKING order="11" place="11" resultid="2677" />
                    <RANKING order="12" place="12" resultid="2093" />
                    <RANKING order="13" place="13" resultid="1811" />
                    <RANKING order="14" place="14" resultid="2551" />
                    <RANKING order="15" place="15" resultid="1516" />
                    <RANKING order="16" place="16" resultid="2080" />
                    <RANKING order="17" place="17" resultid="2548" />
                    <RANKING order="18" place="18" resultid="1486" />
                    <RANKING order="19" place="19" resultid="1844" />
                    <RANKING order="20" place="20" resultid="2659" />
                    <RANKING order="21" place="21" resultid="2043" />
                    <RANKING order="22" place="22" resultid="1791" />
                    <RANKING order="23" place="23" resultid="2202" />
                    <RANKING order="24" place="24" resultid="2521" />
                    <RANKING order="25" place="25" resultid="1209" />
                    <RANKING order="26" place="26" resultid="2475" />
                    <RANKING order="27" place="27" resultid="2483" />
                    <RANKING order="28" place="28" resultid="1587" />
                    <RANKING order="29" place="29" resultid="2529" />
                    <RANKING order="30" place="-1" resultid="1300" />
                    <RANKING order="31" place="-1" resultid="1521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2635" />
                    <RANKING order="2" place="2" resultid="1349" />
                    <RANKING order="3" place="3" resultid="2288" />
                    <RANKING order="4" place="4" resultid="2626" />
                    <RANKING order="5" place="5" resultid="1649" />
                    <RANKING order="6" place="6" resultid="1943" />
                    <RANKING order="7" place="7" resultid="1437" />
                    <RANKING order="8" place="8" resultid="1741" />
                    <RANKING order="9" place="9" resultid="1207" />
                    <RANKING order="10" place="10" resultid="1938" />
                    <RANKING order="11" place="11" resultid="2398" />
                    <RANKING order="12" place="12" resultid="1249" />
                    <RANKING order="13" place="13" resultid="1746" />
                    <RANKING order="14" place="14" resultid="2648" />
                    <RANKING order="15" place="15" resultid="2716" />
                    <RANKING order="16" place="16" resultid="2055" />
                    <RANKING order="17" place="17" resultid="1224" />
                    <RANKING order="18" place="18" resultid="2644" />
                    <RANKING order="19" place="-1" resultid="1536" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3050" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3051" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3052" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3053" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3054" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3055" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="3056" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="3057" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" daytime="14:08" gender="F" number="24" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1152" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1818" />
                    <RANKING order="2" place="2" resultid="2235" />
                    <RANKING order="3" place="3" resultid="2083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="13" agemin="10" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3058" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1155" daytime="14:12" gender="M" number="25" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1156" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2312" />
                    <RANKING order="2" place="2" resultid="2254" />
                    <RANKING order="3" place="3" resultid="1578" />
                    <RANKING order="4" place="4" resultid="2345" />
                    <RANKING order="5" place="5" resultid="1863" />
                    <RANKING order="6" place="6" resultid="1384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="13" agemin="10" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3059" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1159" daytime="14:16" gender="F" number="26" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1160" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2684" />
                    <RANKING order="2" place="2" resultid="2667" />
                    <RANKING order="3" place="3" resultid="1716" />
                    <RANKING order="4" place="4" resultid="1831" />
                    <RANKING order="5" place="5" resultid="2789" />
                    <RANKING order="6" place="6" resultid="2373" />
                    <RANKING order="7" place="7" resultid="2168" />
                    <RANKING order="8" place="8" resultid="2377" />
                    <RANKING order="9" place="9" resultid="2756" />
                    <RANKING order="10" place="10" resultid="1679" />
                    <RANKING order="11" place="11" resultid="1894" />
                    <RANKING order="12" place="12" resultid="2336" />
                    <RANKING order="13" place="13" resultid="2567" />
                    <RANKING order="14" place="14" resultid="2434" />
                    <RANKING order="15" place="15" resultid="2706" />
                    <RANKING order="16" place="16" resultid="1607" />
                    <RANKING order="17" place="17" resultid="2072" />
                    <RANKING order="18" place="18" resultid="1615" />
                    <RANKING order="19" place="19" resultid="1952" />
                    <RANKING order="20" place="20" resultid="1479" />
                    <RANKING order="21" place="21" resultid="1910" />
                    <RANKING order="22" place="22" resultid="2496" />
                    <RANKING order="23" place="23" resultid="2946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1716" />
                    <RANKING order="2" place="2" resultid="2373" />
                    <RANKING order="3" place="3" resultid="2168" />
                    <RANKING order="4" place="4" resultid="2377" />
                    <RANKING order="5" place="5" resultid="2756" />
                    <RANKING order="6" place="6" resultid="1679" />
                    <RANKING order="7" place="7" resultid="1894" />
                    <RANKING order="8" place="8" resultid="2706" />
                    <RANKING order="9" place="9" resultid="2072" />
                    <RANKING order="10" place="10" resultid="1479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2567" />
                    <RANKING order="2" place="2" resultid="1607" />
                    <RANKING order="3" place="3" resultid="1615" />
                    <RANKING order="4" place="4" resultid="1952" />
                    <RANKING order="5" place="5" resultid="1910" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3060" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3061" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3062" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1163" daytime="14:24" gender="M" number="27" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1164" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2730" />
                    <RANKING order="2" place="2" resultid="2795" />
                    <RANKING order="3" place="3" resultid="2595" />
                    <RANKING order="4" place="4" resultid="1279" />
                    <RANKING order="5" place="5" resultid="2779" />
                    <RANKING order="6" place="6" resultid="1508" />
                    <RANKING order="7" place="7" resultid="2743" />
                    <RANKING order="8" place="8" resultid="1238" />
                    <RANKING order="9" place="9" resultid="2552" />
                    <RANKING order="10" place="10" resultid="1767" />
                    <RANKING order="11" place="11" resultid="1517" />
                    <RANKING order="12" place="12" resultid="2387" />
                    <RANKING order="13" place="13" resultid="2660" />
                    <RANKING order="14" place="14" resultid="2308" />
                    <RANKING order="15" place="15" resultid="1835" />
                    <RANKING order="16" place="16" resultid="1526" />
                    <RANKING order="17" place="17" resultid="1847" />
                    <RANKING order="18" place="18" resultid="1201" />
                    <RANKING order="19" place="19" resultid="1588" />
                    <RANKING order="20" place="20" resultid="1998" />
                    <RANKING order="21" place="21" resultid="1583" />
                    <RANKING order="22" place="22" resultid="2580" />
                    <RANKING order="23" place="23" resultid="2586" />
                    <RANKING order="24" place="24" resultid="2562" />
                    <RANKING order="25" place="25" resultid="2283" />
                    <RANKING order="26" place="26" resultid="1732" />
                    <RANKING order="27" place="-1" resultid="1378" />
                    <RANKING order="28" place="-1" resultid="2424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1279" />
                    <RANKING order="2" place="2" resultid="1238" />
                    <RANKING order="3" place="3" resultid="2552" />
                    <RANKING order="4" place="4" resultid="1767" />
                    <RANKING order="5" place="5" resultid="1517" />
                    <RANKING order="6" place="6" resultid="2387" />
                    <RANKING order="7" place="7" resultid="2660" />
                    <RANKING order="8" place="8" resultid="2308" />
                    <RANKING order="9" place="9" resultid="1526" />
                    <RANKING order="10" place="10" resultid="1847" />
                    <RANKING order="11" place="11" resultid="1588" />
                    <RANKING order="12" place="-1" resultid="1378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1201" />
                    <RANKING order="2" place="2" resultid="1998" />
                    <RANKING order="3" place="3" resultid="1583" />
                    <RANKING order="4" place="4" resultid="2283" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3063" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3064" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3065" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1167" daytime="14:32" gender="F" number="28" order="29" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1168" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2685" />
                    <RANKING order="2" place="2" resultid="2240" />
                    <RANKING order="3" place="3" resultid="2792" />
                    <RANKING order="4" place="4" resultid="2180" />
                    <RANKING order="5" place="5" resultid="2265" />
                    <RANKING order="6" place="6" resultid="2381" />
                    <RANKING order="7" place="7" resultid="2354" />
                    <RANKING order="8" place="8" resultid="2084" />
                    <RANKING order="9" place="9" resultid="2278" />
                    <RANKING order="10" place="10" resultid="2325" />
                    <RANKING order="11" place="11" resultid="2341" />
                    <RANKING order="12" place="12" resultid="2214" />
                    <RANKING order="13" place="13" resultid="1780" />
                    <RANKING order="14" place="14" resultid="2192" />
                    <RANKING order="15" place="15" resultid="1977" />
                    <RANKING order="16" place="16" resultid="2333" />
                    <RANKING order="17" place="17" resultid="1611" />
                    <RANKING order="18" place="18" resultid="2443" />
                    <RANKING order="19" place="19" resultid="1623" />
                    <RANKING order="20" place="20" resultid="2623" />
                    <RANKING order="21" place="21" resultid="3083" />
                    <RANKING order="22" place="22" resultid="1927" />
                    <RANKING order="23" place="23" resultid="1229" />
                    <RANKING order="24" place="24" resultid="1957" />
                    <RANKING order="25" place="-1" resultid="1455" />
                    <RANKING order="26" place="-1" resultid="1546" />
                    <RANKING order="27" place="-1" resultid="1628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2240" />
                    <RANKING order="2" place="2" resultid="2792" />
                    <RANKING order="3" place="3" resultid="2265" />
                    <RANKING order="4" place="4" resultid="2381" />
                    <RANKING order="5" place="5" resultid="2354" />
                    <RANKING order="6" place="6" resultid="2084" />
                    <RANKING order="7" place="7" resultid="2278" />
                    <RANKING order="8" place="8" resultid="2325" />
                    <RANKING order="9" place="9" resultid="2341" />
                    <RANKING order="10" place="10" resultid="2214" />
                    <RANKING order="11" place="11" resultid="2192" />
                    <RANKING order="12" place="12" resultid="2333" />
                    <RANKING order="13" place="13" resultid="2443" />
                    <RANKING order="14" place="14" resultid="1623" />
                    <RANKING order="15" place="-1" resultid="1455" />
                    <RANKING order="16" place="-1" resultid="1546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1780" />
                    <RANKING order="2" place="2" resultid="1977" />
                    <RANKING order="3" place="3" resultid="1611" />
                    <RANKING order="4" place="4" resultid="2623" />
                    <RANKING order="5" place="5" resultid="3083" />
                    <RANKING order="6" place="6" resultid="1927" />
                    <RANKING order="7" place="7" resultid="1229" />
                    <RANKING order="8" place="8" resultid="1957" />
                    <RANKING order="9" place="-1" resultid="1628" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3066" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3067" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3068" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1171" daytime="14:44" gender="M" number="29" order="30" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1172" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                    <RANKING order="2" place="2" resultid="2804" />
                    <RANKING order="3" place="3" resultid="1727" />
                    <RANKING order="4" place="4" resultid="2259" />
                    <RANKING order="5" place="5" resultid="2183" />
                    <RANKING order="6" place="6" resultid="2296" />
                    <RANKING order="7" place="7" resultid="1661" />
                    <RANKING order="8" place="8" resultid="1879" />
                    <RANKING order="9" place="9" resultid="1987" />
                    <RANKING order="10" place="10" resultid="1752" />
                    <RANKING order="11" place="11" resultid="1338" />
                    <RANKING order="12" place="12" resultid="1640" />
                    <RANKING order="13" place="13" resultid="1447" />
                    <RANKING order="14" place="14" resultid="1504" />
                    <RANKING order="15" place="15" resultid="2661" />
                    <RANKING order="16" place="16" resultid="1982" />
                    <RANKING order="17" place="17" resultid="2250" />
                    <RANKING order="18" place="18" resultid="1991" />
                    <RANKING order="19" place="19" resultid="2206" />
                    <RANKING order="20" place="20" resultid="1742" />
                    <RANKING order="21" place="21" resultid="2399" />
                    <RANKING order="22" place="22" resultid="1650" />
                    <RANKING order="23" place="23" resultid="1273" />
                    <RANKING order="24" place="24" resultid="1737" />
                    <RANKING order="25" place="25" resultid="1747" />
                    <RANKING order="26" place="26" resultid="2627" />
                    <RANKING order="27" place="-1" resultid="2649" />
                    <RANKING order="28" place="-1" resultid="1785" />
                    <RANKING order="29" place="-1" resultid="1807" />
                    <RANKING order="30" place="-1" resultid="1851" />
                    <RANKING order="31" place="-1" resultid="2425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                    <RANKING order="2" place="2" resultid="2804" />
                    <RANKING order="3" place="3" resultid="2259" />
                    <RANKING order="4" place="4" resultid="2183" />
                    <RANKING order="5" place="5" resultid="1661" />
                    <RANKING order="6" place="6" resultid="1879" />
                    <RANKING order="7" place="7" resultid="1987" />
                    <RANKING order="8" place="8" resultid="1640" />
                    <RANKING order="9" place="9" resultid="2661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2250" />
                    <RANKING order="2" place="2" resultid="1991" />
                    <RANKING order="3" place="3" resultid="2206" />
                    <RANKING order="4" place="4" resultid="1742" />
                    <RANKING order="5" place="5" resultid="2399" />
                    <RANKING order="6" place="6" resultid="1650" />
                    <RANKING order="7" place="7" resultid="1747" />
                    <RANKING order="8" place="8" resultid="2627" />
                    <RANKING order="9" place="-1" resultid="2649" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3069" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3070" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3071" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3072" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1175" daytime="15:00" gender="F" number="30" order="31" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1176" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1860" />
                    <RANKING order="2" place="2" resultid="1441" />
                    <RANKING order="3" place="3" resultid="1392" />
                    <RANKING order="4" place="4" resultid="1598" />
                    <RANKING order="5" place="5" resultid="1965" />
                    <RANKING order="6" place="6" resultid="2132" />
                    <RANKING order="7" place="7" resultid="1361" />
                    <RANKING order="8" place="8" resultid="1242" />
                    <RANKING order="9" place="9" resultid="1387" />
                    <RANKING order="10" place="10" resultid="1856" />
                    <RANKING order="11" place="11" resultid="1358" />
                    <RANKING order="12" place="-1" resultid="2304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1441" />
                    <RANKING order="2" place="2" resultid="1392" />
                    <RANKING order="3" place="3" resultid="1598" />
                    <RANKING order="4" place="4" resultid="1965" />
                    <RANKING order="5" place="-1" resultid="2304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1361" />
                    <RANKING order="2" place="2" resultid="1242" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3073" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3074" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1179" daytime="15:14" gender="M" number="31" order="32" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1180" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2570" />
                    <RANKING order="2" place="2" resultid="2769" />
                    <RANKING order="3" place="3" resultid="1868" />
                    <RANKING order="4" place="4" resultid="2573" />
                    <RANKING order="5" place="5" resultid="1496" />
                    <RANKING order="6" place="6" resultid="1245" />
                    <RANKING order="7" place="7" resultid="2537" />
                    <RANKING order="8" place="8" resultid="2120" />
                    <RANKING order="9" place="9" resultid="2616" />
                    <RANKING order="10" place="10" resultid="2576" />
                    <RANKING order="11" place="11" resultid="1409" />
                    <RANKING order="12" place="12" resultid="1645" />
                    <RANKING order="13" place="13" resultid="1864" />
                    <RANKING order="14" place="14" resultid="1836" />
                    <RANKING order="15" place="15" resultid="1250" />
                    <RANKING order="16" place="16" resultid="1385" />
                    <RANKING order="17" place="17" resultid="1324" />
                    <RANKING order="18" place="18" resultid="2556" />
                    <RANKING order="19" place="19" resultid="1304" />
                    <RANKING order="20" place="-1" resultid="1872" />
                    <RANKING order="21" place="-1" resultid="2125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="16" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1245" />
                    <RANKING order="2" place="2" resultid="2537" />
                    <RANKING order="3" place="3" resultid="2616" />
                    <RANKING order="4" place="4" resultid="2576" />
                    <RANKING order="5" place="5" resultid="1409" />
                    <RANKING order="6" place="6" resultid="1645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="13" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2120" />
                    <RANKING order="2" place="2" resultid="1250" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3075" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3076" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3077" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" daytime="15:32" gender="X" number="32" order="33" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1184" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2186" />
                    <RANKING order="2" place="2" resultid="1886" />
                    <RANKING order="3" place="3" resultid="2187" />
                    <RANKING order="4" place="4" resultid="2360" />
                    <RANKING order="5" place="5" resultid="2361" />
                    <RANKING order="6" place="6" resultid="1601" />
                    <RANKING order="7" place="7" resultid="1887" />
                    <RANKING order="8" place="8" resultid="2362" />
                    <RANKING order="9" place="9" resultid="1655" />
                    <RANKING order="10" place="10" resultid="1959" />
                    <RANKING order="11" place="11" resultid="1960" />
                    <RANKING order="12" place="-1" resultid="2359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="16" agemin="14" />
                <AGEGROUP agegroupid="1186" agemax="13" agemin="10" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3078" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3079" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="06401" nation="POL" region="01" clubid="1339" name="KS &quot;Swimmers Centrum Ślęza&quot;">
          <ATHLETES>
            <ATHLETE firstname="Radosław" lastname="Stefurak" birthdate="1974-09-07" gender="M" nation="POL" license="506401700019" swrid="4429483" athleteid="1350">
              <RESULTS>
                <RESULT eventid="1083" reactiontime="+93" status="DNF" swimtime="00:00:00.00" resultid="1351" heatid="2974" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                    <SPLIT distance="100" swimtime="00:01:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="257" reactiontime="+101" swimtime="00:01:29.35" resultid="1352" heatid="3007" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="269" reactiontime="+97" swimtime="00:00:40.18" resultid="1353" heatid="3054" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Wolny" birthdate="1960-03-21" gender="M" nation="POL" license="506401700021" swrid="4183808" athleteid="1354">
              <RESULTS>
                <RESULT eventid="1099" points="349" reactiontime="+69" swimtime="00:00:34.08" resultid="1355" heatid="2990" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Wolny" birthdate="2011-04-18" gender="M" nation="POL" license="106401700018" swrid="5461258" athleteid="1343">
              <RESULTS>
                <RESULT eventid="1075" points="153" swimtime="00:00:39.07" resultid="1344" heatid="2960" lane="8" />
                <RESULT eventid="1099" points="167" reactiontime="+57" swimtime="00:00:43.58" resultid="1345" heatid="2989" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Burandt" birthdate="2011-03-19" gender="F" nation="POL" license="106401600010" swrid="5217597" athleteid="1340">
              <RESULTS>
                <RESULT eventid="1071" points="253" reactiontime="+90" swimtime="00:00:37.41" resultid="1341" heatid="2951" lane="8" />
                <RESULT eventid="1119" points="139" reactiontime="+89" swimtime="00:00:47.10" resultid="1342" heatid="3013" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pola" lastname="Pietryk" birthdate="2008-09-26" gender="F" nation="POL" license="106401600002" swrid="5354927" athleteid="1359">
              <RESULTS>
                <RESULT eventid="1103" points="400" reactiontime="+85" swimtime="00:02:33.30" resultid="1360" heatid="2996" lane="0" entrytime="00:02:35.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:13.88" />
                    <SPLIT distance="150" swimtime="00:01:54.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="370" reactiontime="+86" swimtime="00:05:29.26" resultid="1361" heatid="3074" lane="1" entrytime="00:05:25.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:01:17.34" />
                    <SPLIT distance="150" swimtime="00:01:58.56" />
                    <SPLIT distance="200" swimtime="00:02:40.78" />
                    <SPLIT distance="250" swimtime="00:03:24.54" />
                    <SPLIT distance="300" swimtime="00:04:07.76" />
                    <SPLIT distance="350" swimtime="00:04:50.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julian" lastname="Stefurak" birthdate="2008-05-02" gender="M" nation="POL" license="106401700004" swrid="5311183" athleteid="1346">
              <RESULTS>
                <RESULT eventid="1083" points="267" reactiontime="+75" swimtime="00:03:15.82" resultid="1347" heatid="2975" lane="4" entrytime="00:03:07.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                    <SPLIT distance="100" swimtime="00:01:34.07" />
                    <SPLIT distance="150" swimtime="00:02:25.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="249" reactiontime="+67" swimtime="00:01:30.33" resultid="1348" heatid="3008" lane="3" entrytime="00:01:26.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="295" reactiontime="+65" swimtime="00:00:38.98" resultid="1349" heatid="3055" lane="5" entrytime="00:00:38.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Burandt" birthdate="1972-12-15" gender="F" nation="POL" license="506401600020" athleteid="1356">
              <RESULTS>
                <RESULT eventid="1103" points="216" reactiontime="+115" swimtime="00:03:08.19" resultid="1357" heatid="2995" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                    <SPLIT distance="100" swimtime="00:01:25.26" />
                    <SPLIT distance="150" swimtime="00:02:16.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="207" swimtime="00:06:39.44" resultid="1358" heatid="3073" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                    <SPLIT distance="100" swimtime="00:01:29.17" />
                    <SPLIT distance="150" swimtime="00:02:18.59" />
                    <SPLIT distance="200" swimtime="00:03:08.99" />
                    <SPLIT distance="250" swimtime="00:04:00.86" />
                    <SPLIT distance="300" swimtime="00:04:53.71" />
                    <SPLIT distance="350" swimtime="00:05:46.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02915" nation="POL" region="15" clubid="2455" name="UKS 3-Wodnik Wolsztyn">
          <ATHLETES>
            <ATHLETE firstname="Magdalena" lastname="Dechnik" birthdate="2008-09-26" gender="F" nation="POL" license="102915600077" swrid="5254262" athleteid="2456">
              <RESULTS>
                <RESULT eventid="1071" points="289" reactiontime="+103" swimtime="00:00:35.79" resultid="2457" heatid="2952" lane="7" />
                <RESULT eventid="1135" points="272" reactiontime="+88" swimtime="00:01:19.78" resultid="2458" heatid="3029" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="295" reactiontime="+91" swimtime="00:00:44.13" resultid="2459" heatid="3045" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Weiss" birthdate="2008-05-27" gender="F" nation="POL" license="102915600093" swrid="5342869" athleteid="2460">
              <RESULTS>
                <RESULT eventid="1071" points="225" reactiontime="+90" swimtime="00:00:38.89" resultid="2461" heatid="2951" lane="4" />
                <RESULT eventid="1095" points="198" reactiontime="+64" swimtime="00:00:46.23" resultid="2462" heatid="2985" lane="5" entrytime="00:00:46.49" entrycourse="LCM" />
                <RESULT eventid="1119" points="118" reactiontime="+75" swimtime="00:00:49.68" resultid="2463" heatid="3013" lane="5" entrytime="00:00:48.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Sławiński" birthdate="2006-10-16" gender="M" nation="POL" license="102915700069" swrid="4838415" athleteid="2476">
              <RESULTS>
                <RESULT eventid="1075" points="271" reactiontime="+89" swimtime="00:00:32.29" resultid="2477" heatid="2961" lane="3" />
                <RESULT eventid="1123" points="221" reactiontime="+82" swimtime="00:00:36.79" resultid="2478" heatid="3019" lane="6" />
                <RESULT eventid="1139" points="262" reactiontime="+83" swimtime="00:01:13.25" resultid="2479" heatid="3037" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymon" lastname="Grabczyński" birthdate="2007-02-16" gender="M" nation="POL" license="102915700107" swrid="5342857" athleteid="2472">
              <RESULTS>
                <RESULT eventid="1075" points="326" reactiontime="+74" swimtime="00:00:30.38" resultid="2473" heatid="2967" lane="7" entrytime="00:00:29.91" entrycourse="LCM" />
                <RESULT eventid="1123" points="213" reactiontime="+81" swimtime="00:00:37.25" resultid="2474" heatid="3019" lane="9" />
                <RESULT eventid="1147" points="242" reactiontime="+78" swimtime="00:00:41.61" resultid="2475" heatid="3051" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Kasperowicz" birthdate="2008-04-06" gender="F" nation="POL" license="102915600083" swrid="5254260" athleteid="2484">
              <RESULTS>
                <RESULT eventid="1079" points="325" reactiontime="+92" swimtime="00:03:22.17" resultid="2485" heatid="2973" lane="9" entrytime="00:03:29.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                    <SPLIT distance="100" swimtime="00:01:35.61" />
                    <SPLIT distance="150" swimtime="00:02:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="349" reactiontime="+91" swimtime="00:01:31.05" resultid="2486" heatid="3004" lane="1" entrytime="00:01:31.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="392" reactiontime="+84" swimtime="00:00:40.16" resultid="2487" heatid="3048" lane="0" entrytime="00:00:40.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Wojtkowiak" birthdate="2007-12-22" gender="M" nation="POL" license="102915700082" swrid="5254258" athleteid="2468">
              <RESULTS>
                <RESULT eventid="1075" points="361" reactiontime="+83" swimtime="00:00:29.35" resultid="2469" heatid="2966" lane="4" entrytime="00:00:30.59" entrycourse="LCM" />
                <RESULT eventid="1099" points="322" reactiontime="+72" swimtime="00:00:34.98" resultid="2470" heatid="2988" lane="4" />
                <RESULT eventid="1123" points="251" reactiontime="+90" swimtime="00:00:35.30" resultid="2471" heatid="3018" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Tomys" birthdate="2005-08-31" gender="M" nation="POL" license="102915700055" swrid="5162122" athleteid="2464">
              <RESULTS>
                <RESULT eventid="1075" points="366" reactiontime="+82" swimtime="00:00:29.22" resultid="2465" heatid="2968" lane="8" entrytime="00:00:28.64" entrycourse="LCM" />
                <RESULT eventid="1123" points="304" reactiontime="+74" swimtime="00:00:33.12" resultid="2466" heatid="3020" lane="0" />
                <RESULT eventid="1139" points="394" reactiontime="+74" swimtime="00:01:03.98" resultid="2467" heatid="3039" lane="3" entrytime="00:01:03.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Wieczorek" birthdate="2007-02-25" gender="M" nation="POL" license="102915700088" swrid="5342872" athleteid="2480">
              <RESULTS>
                <RESULT eventid="1075" points="238" reactiontime="+104" swimtime="00:00:33.72" resultid="2481" heatid="2964" lane="9" />
                <RESULT eventid="1115" points="240" reactiontime="+91" swimtime="00:01:31.42" resultid="2482" heatid="3008" lane="7" entrytime="00:01:32.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="238" swimtime="00:00:41.87" resultid="2483" heatid="3055" lane="2" entrytime="00:00:41.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05201" nation="POL" region="01" clubid="1380" name="KS JUST SWIM Jelenia Góra">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Lara" birthdate="1985-06-16" gender="F" nation="POL" license="505201600088" swrid="5435203" athleteid="1386">
              <RESULTS>
                <RESULT eventid="1175" points="234" reactiontime="+100" swimtime="00:06:23.47" resultid="1387" heatid="3073" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:01:27.97" />
                    <SPLIT distance="150" swimtime="00:02:17.17" />
                    <SPLIT distance="200" swimtime="00:03:05.97" />
                    <SPLIT distance="250" swimtime="00:03:56.21" />
                    <SPLIT distance="300" swimtime="00:04:44.84" />
                    <SPLIT distance="350" swimtime="00:05:35.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Lipka" birthdate="1958-06-05" gender="M" nation="POL" license="505201700087" swrid="5435204" athleteid="1381">
              <RESULTS>
                <RESULT eventid="1091" points="111" reactiontime="+104" swimtime="00:01:42.81" resultid="1382" heatid="2980" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="153" reactiontime="+106" swimtime="00:03:10.44" resultid="1383" heatid="2999" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:32.94" />
                    <SPLIT distance="150" swimtime="00:02:23.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="102" reactiontime="+93" swimtime="00:03:56.93" resultid="1384" heatid="3059" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.07" />
                    <SPLIT distance="100" swimtime="00:01:53.10" />
                    <SPLIT distance="150" swimtime="00:02:53.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="165" reactiontime="+94" swimtime="00:06:40.76" resultid="1385" heatid="3076" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.43" />
                    <SPLIT distance="100" swimtime="00:01:36.50" />
                    <SPLIT distance="150" swimtime="00:02:27.96" />
                    <SPLIT distance="200" swimtime="00:03:19.82" />
                    <SPLIT distance="250" swimtime="00:04:11.97" />
                    <SPLIT distance="300" swimtime="00:05:05.07" />
                    <SPLIT distance="350" swimtime="00:05:54.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00101" nation="POL" region="01" clubid="2146" name="MKS Juvenia Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Maja" lastname="Malaczewska" birthdate="2005-07-05" gender="F" nation="POL" license="100101601336" swrid="5088657" athleteid="2166">
              <RESULTS>
                <RESULT eventid="1103" points="533" reactiontime="+69" swimtime="00:02:19.30" resultid="2167" heatid="2996" lane="4" entrytime="00:02:20.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                    <SPLIT distance="100" swimtime="00:01:06.76" />
                    <SPLIT distance="150" swimtime="00:01:43.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="550" reactiontime="+69" swimtime="00:01:10.26" resultid="2168" heatid="3062" lane="7" entrytime="00:01:09.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Maciuszek" birthdate="2004-05-11" gender="F" nation="POL" license="100101601407" swrid="4858842" athleteid="2147">
              <RESULTS>
                <RESULT eventid="1071" points="643" reactiontime="+67" swimtime="00:00:27.41" resultid="2148" heatid="2959" lane="4" entrytime="00:00:27.19" entrycourse="LCM" />
                <RESULT eventid="1095" points="694" reactiontime="+55" swimtime="00:00:30.47" resultid="2149" heatid="2987" lane="5" entrytime="00:00:30.56" entrycourse="LCM" />
                <RESULT eventid="1119" points="585" reactiontime="+71" swimtime="00:00:29.20" resultid="2150" heatid="3016" lane="3" entrytime="00:00:29.43" entrycourse="LCM" />
                <RESULT eventid="1143" points="570" reactiontime="+72" swimtime="00:00:35.45" resultid="2151" heatid="3046" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Sarnowicz" birthdate="2004-03-01" gender="M" nation="POL" license="100101701073" swrid="5118745" athleteid="2175">
              <RESULTS>
                <RESULT eventid="1123" points="478" reactiontime="+68" swimtime="00:00:28.48" resultid="2176" heatid="3018" lane="0" />
                <RESULT eventid="1139" points="518" reactiontime="+68" swimtime="00:00:58.41" resultid="2177" heatid="3035" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Strużyk" birthdate="2004-06-27" gender="F" nation="POL" license="100101601049" swrid="5072852" athleteid="2178">
              <RESULTS>
                <RESULT eventid="1135" points="557" reactiontime="+80" swimtime="00:01:02.83" resultid="2179" heatid="3030" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="545" reactiontime="+75" swimtime="00:02:34.34" resultid="2180" heatid="3068" lane="3" entrytime="00:02:33.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:56.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alex" lastname="Rytkowski" birthdate="2005-03-21" gender="M" nation="POL" license="100101701227" swrid="5113513" athleteid="2169">
              <RESULTS>
                <RESULT eventid="1115" points="531" reactiontime="+75" swimtime="00:01:10.20" resultid="2170" heatid="3009" lane="4" entrytime="00:01:10.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="539" reactiontime="+67" swimtime="00:00:31.88" resultid="2171" heatid="3057" lane="1" entrytime="00:00:31.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Malwina" lastname="Malaczewska" birthdate="2005-07-05" gender="F" nation="POL" license="100101601337" swrid="5088658" athleteid="2158">
              <RESULTS>
                <RESULT eventid="1071" points="636" reactiontime="+58" swimtime="00:00:27.51" resultid="2159" heatid="2959" lane="5" entrytime="00:00:27.22" entrycourse="LCM" />
                <RESULT eventid="1135" points="635" reactiontime="+69" swimtime="00:01:00.16" resultid="2160" heatid="3034" lane="6" entrytime="00:01:00.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Durlik" birthdate="2005-04-30" gender="M" nation="POL" license="100101701335" swrid="5118820" athleteid="2172">
              <RESULTS>
                <RESULT eventid="1123" points="539" reactiontime="+57" swimtime="00:00:27.36" resultid="2173" heatid="3023" lane="5" entrytime="00:00:27.45" entrycourse="LCM" />
                <RESULT eventid="1139" points="533" reactiontime="+70" swimtime="00:00:57.84" resultid="2174" heatid="3041" lane="7" entrytime="00:00:58.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Kramkowska" birthdate="2004-09-29" gender="F" nation="POL" license="100101601287" swrid="4990815" athleteid="2161">
              <RESULTS>
                <RESULT eventid="1071" points="562" reactiontime="+75" swimtime="00:00:28.67" resultid="2162" heatid="2959" lane="8" entrytime="00:00:28.25" entrycourse="LCM" />
                <RESULT eventid="1087" points="498" reactiontime="+74" swimtime="00:01:09.95" resultid="2163" heatid="2978" lane="3" entrytime="00:01:08.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="546" reactiontime="+77" swimtime="00:01:03.26" resultid="2164" heatid="3034" lane="8" entrytime="00:01:01.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Wierzbicki" birthdate="2005-06-25" gender="M" nation="POL" license="100101701334" swrid="5147678" athleteid="2181">
              <RESULTS>
                <RESULT eventid="1139" points="555" reactiontime="+66" swimtime="00:00:57.05" resultid="2182" heatid="3042" lane="0" entrytime="00:00:57.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="516" reactiontime="+68" swimtime="00:02:22.06" resultid="2183" heatid="3072" lane="6" entrytime="00:02:20.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                    <SPLIT distance="100" swimtime="00:01:05.58" />
                    <SPLIT distance="150" swimtime="00:01:49.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iga" lastname="Maślej" birthdate="2003-05-15" gender="F" nation="POL" license="100101601020" swrid="5043142" athleteid="2152">
              <RESULTS>
                <RESULT eventid="1071" points="506" reactiontime="+75" swimtime="00:00:29.69" resultid="2153" heatid="2958" lane="9" entrytime="00:00:29.27" entrycourse="LCM" />
                <RESULT eventid="1087" points="505" reactiontime="+73" swimtime="00:01:09.65" resultid="2154" heatid="2978" lane="6" entrytime="00:01:09.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="556" reactiontime="+70" swimtime="00:02:17.33" resultid="2155" heatid="2997" lane="7" entrytime="00:02:16.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:06.58" />
                    <SPLIT distance="150" swimtime="00:01:42.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="461" swimtime="00:00:31.62" resultid="2156" heatid="3015" lane="2" entrytime="00:00:31.36" entrycourse="LCM" />
                <RESULT eventid="1135" points="537" swimtime="00:01:03.58" resultid="2157" heatid="3033" lane="2" entrytime="00:01:03.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+68" swimtime="00:01:47.20" resultid="2184" heatid="2947" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.83" />
                    <SPLIT distance="100" swimtime="00:00:53.07" />
                    <SPLIT distance="150" swimtime="00:01:20.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2172" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2166" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="2158" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="2181" number="4" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1183" reactiontime="+64" swimtime="00:01:57.42" resultid="2186" heatid="3078" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:02.89" />
                    <SPLIT distance="150" swimtime="00:01:29.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2178" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2175" number="2" reactiontime="-1" />
                    <RELAYPOSITION athleteid="2172" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="2161" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1059" swimtime="00:01:48.93" resultid="2185" heatid="2947" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                    <SPLIT distance="100" swimtime="00:00:53.88" />
                    <SPLIT distance="150" swimtime="00:01:22.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2169" number="1" />
                    <RELAYPOSITION athleteid="2178" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2152" number="3" />
                    <RELAYPOSITION athleteid="2175" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1183" reactiontime="+64" swimtime="00:01:59.10" resultid="2187" heatid="3079" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:05.81" />
                    <SPLIT distance="150" swimtime="00:01:33.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2166" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2158" number="2" />
                    <RELAYPOSITION athleteid="2181" number="3" reactiontime="+1" />
                    <RELAYPOSITION athleteid="2169" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00315" nation="POL" region="15" clubid="2017" name="MKP Astromal-Leszno">
          <ATHLETES>
            <ATHLETE firstname="Oliwia" lastname="Juszkiewicz" birthdate="2007-12-06" gender="F" nation="POL" license="100315600389" swrid="5298518" athleteid="2068">
              <RESULTS>
                <RESULT eventid="1079" points="478" reactiontime="+55" swimtime="00:02:57.87" resultid="2069" heatid="2973" lane="2" entrytime="00:03:02.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:01:24.06" />
                    <SPLIT distance="150" swimtime="00:02:10.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="459" reactiontime="+81" swimtime="00:01:23.12" resultid="2070" heatid="3005" lane="8" entrytime="00:01:21.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="497" reactiontime="+71" swimtime="00:00:37.10" resultid="2071" heatid="3049" lane="0" entrytime="00:00:36.80" entrycourse="LCM" />
                <RESULT eventid="1159" points="361" reactiontime="+71" swimtime="00:01:20.83" resultid="2072" heatid="3060" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Błazik" birthdate="2008-04-29" gender="F" nation="POL" license="100315600382" swrid="5311261" athleteid="2022">
              <RESULTS>
                <RESULT eventid="1071" points="306" reactiontime="+74" swimtime="00:00:35.11" resultid="2023" heatid="2953" lane="1" />
                <RESULT eventid="1095" points="257" reactiontime="+84" swimtime="00:00:42.42" resultid="2024" heatid="2986" lane="9" entrytime="00:00:41.88" entrycourse="LCM" />
                <RESULT eventid="1135" points="291" swimtime="00:01:18.00" resultid="2025" heatid="3030" lane="2" entrytime="00:01:22.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Staniewski" birthdate="2006-09-07" gender="M" nation="POL" license="100315700367" swrid="4952524" athleteid="2073">
              <RESULTS>
                <RESULT eventid="1083" points="376" reactiontime="+72" swimtime="00:02:54.71" resultid="2074" heatid="2976" lane="0" entrytime="00:02:55.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:23.31" />
                    <SPLIT distance="150" swimtime="00:02:09.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="398" reactiontime="+85" swimtime="00:01:17.27" resultid="2075" heatid="3007" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Uzarowski" birthdate="2006-07-20" gender="M" nation="POL" license="100315700370" swrid="4951994" athleteid="2033">
              <RESULTS>
                <RESULT eventid="1075" points="276" reactiontime="+82" swimtime="00:00:32.10" resultid="2034" heatid="2966" lane="8" entrytime="00:00:32.21" entrycourse="LCM" />
                <RESULT eventid="1107" points="262" reactiontime="+82" swimtime="00:02:39.35" resultid="2035" heatid="3000" lane="8" entrytime="00:02:41.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:17.24" />
                    <SPLIT distance="150" swimtime="00:01:59.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="270" reactiontime="+70" swimtime="00:01:12.54" resultid="2036" heatid="3038" lane="6" entrytime="00:01:12.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Szarszewski" birthdate="2007-10-01" gender="M" nation="POL" license="100315700401" swrid="5298516" athleteid="2076">
              <RESULTS>
                <RESULT eventid="1083" points="389" reactiontime="+73" swimtime="00:02:52.64" resultid="2077" heatid="2975" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                    <SPLIT distance="100" swimtime="00:01:24.85" />
                    <SPLIT distance="150" swimtime="00:02:09.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1091" points="284" reactiontime="+88" swimtime="00:01:15.27" resultid="2078" heatid="2981" lane="7" entrytime="00:01:15.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="360" reactiontime="+74" swimtime="00:01:19.89" resultid="2079" heatid="3009" lane="9" entrytime="00:01:18.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="365" reactiontime="+70" swimtime="00:00:36.30" resultid="2080" heatid="3052" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Budzeń" birthdate="2007-07-18" gender="F" nation="POL" license="100315600384" swrid="5298519" athleteid="2081">
              <RESULTS>
                <RESULT eventid="1087" points="473" swimtime="00:01:11.20" resultid="2082" heatid="2978" lane="2" entrytime="00:01:12.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="445" reactiontime="+80" swimtime="00:02:39.50" resultid="2083" heatid="3058" lane="3" entrytime="00:02:47.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:14.23" />
                    <SPLIT distance="150" swimtime="00:01:56.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="477" reactiontime="+87" swimtime="00:02:41.37" resultid="2084" heatid="3067" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                    <SPLIT distance="100" swimtime="00:01:20.33" />
                    <SPLIT distance="150" swimtime="00:02:06.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Kozłowski" birthdate="2007-10-11" gender="M" nation="POL" license="100315700390" swrid="5311255" athleteid="2044">
              <RESULTS>
                <RESULT eventid="1075" points="228" reactiontime="+90" swimtime="00:00:34.18" resultid="2045" heatid="2964" lane="2" />
                <RESULT eventid="1099" points="199" reactiontime="+71" swimtime="00:00:41.06" resultid="2046" heatid="2989" lane="6" />
                <RESULT eventid="1139" points="242" reactiontime="+89" swimtime="00:01:15.19" resultid="2047" heatid="3036" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Janiak" birthdate="2007-03-28" gender="M" nation="POL" license="100315700358" swrid="4951953" athleteid="2091">
              <RESULTS>
                <RESULT eventid="1115" points="417" reactiontime="+62" swimtime="00:01:16.11" resultid="2092" heatid="3009" lane="0" entrytime="00:01:15.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="426" reactiontime="+72" swimtime="00:00:34.47" resultid="2093" heatid="3056" lane="7" entrytime="00:00:34.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Jakubiak" birthdate="2005-07-25" gender="M" nation="POL" license="100315700329" swrid="5153463" athleteid="2056">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="2057" heatid="2967" lane="4" entrytime="00:00:29.14" entrycourse="LCM" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="2058" heatid="3039" lane="4" entrytime="00:01:03.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymoteusz" lastname="Wołowicz" birthdate="2006-05-20" gender="M" nation="POL" license="100315700372" swrid="5202110" athleteid="2085">
              <RESULTS>
                <RESULT eventid="1091" points="491" reactiontime="+70" swimtime="00:01:02.72" resultid="2086" heatid="2982" lane="1" entrytime="00:01:01.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="524" reactiontime="+72" swimtime="00:00:27.61" resultid="2087" heatid="3023" lane="6" entrytime="00:00:27.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Krawczyk" birthdate="2007-06-19" gender="F" nation="POL" license="100315600381" swrid="5204394" athleteid="2018">
              <RESULTS>
                <RESULT eventid="1071" points="421" reactiontime="+79" swimtime="00:00:31.57" resultid="2019" heatid="2951" lane="5" />
                <RESULT eventid="1095" points="383" reactiontime="+79" swimtime="00:00:37.12" resultid="2020" heatid="2986" lane="1" entrytime="00:00:38.23" entrycourse="LCM" />
                <RESULT eventid="1143" points="393" reactiontime="+79" swimtime="00:00:40.12" resultid="2021" heatid="3046" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tobiasz" lastname="Walkowski" birthdate="2006-11-25" gender="M" nation="POL" license="100315700371" swrid="4951851" athleteid="2037">
              <RESULTS>
                <RESULT eventid="1075" points="331" reactiontime="+95" swimtime="00:00:30.21" resultid="2038" heatid="2963" lane="7" />
                <RESULT eventid="1139" points="360" reactiontime="+73" swimtime="00:01:05.91" resultid="2039" heatid="3039" lane="1" entrytime="00:01:05.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Godzisz" birthdate="2006-02-27" gender="M" nation="POL" license="100315700353" swrid="4951850" athleteid="2029">
              <RESULTS>
                <RESULT eventid="1075" points="460" reactiontime="+75" swimtime="00:00:27.08" resultid="2030" heatid="2968" lane="5" entrytime="00:00:27.63" entrycourse="LCM" />
                <RESULT eventid="1107" points="414" reactiontime="+83" swimtime="00:02:16.75" resultid="2031" heatid="3000" lane="6" entrytime="00:02:18.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:05.68" />
                    <SPLIT distance="150" swimtime="00:01:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="490" reactiontime="+71" swimtime="00:00:59.48" resultid="2032" heatid="3041" lane="0" entrytime="00:00:59.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Stawiński" birthdate="2007-12-08" gender="M" nation="POL" license="100315700400" swrid="5298514" athleteid="2040">
              <RESULTS>
                <RESULT eventid="1075" points="339" reactiontime="+77" swimtime="00:00:29.98" resultid="2041" heatid="2967" lane="9" entrytime="00:00:30.19" entrycourse="LCM" />
                <RESULT eventid="1115" points="304" reactiontime="+74" swimtime="00:01:24.54" resultid="2042" heatid="3008" lane="5" entrytime="00:01:25.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="317" reactiontime="+77" swimtime="00:00:38.04" resultid="2043" heatid="3056" lane="9" entrytime="00:00:36.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Grining" birthdate="2006-02-18" gender="M" nation="POL" license="100315700355" swrid="4951946" athleteid="2088">
              <RESULTS>
                <RESULT eventid="1091" points="305" reactiontime="+67" swimtime="00:01:13.53" resultid="2089" heatid="2981" lane="2" entrytime="00:01:11.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="352" reactiontime="+76" swimtime="00:01:06.38" resultid="2090" heatid="3039" lane="7" entrytime="00:01:04.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kinga" lastname="Przybysz" birthdate="2004-11-05" gender="F" nation="POL" license="100315600318" swrid="5114696" athleteid="2026">
              <RESULTS>
                <RESULT eventid="1071" points="498" reactiontime="+87" swimtime="00:00:29.86" resultid="2027" heatid="2953" lane="3" />
                <RESULT eventid="1079" points="464" reactiontime="+83" swimtime="00:02:59.67" resultid="2028" heatid="2973" lane="6" entrytime="00:02:58.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:27.40" />
                    <SPLIT distance="150" swimtime="00:02:13.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Janiak" birthdate="2005-01-21" gender="M" nation="POL" license="100315700307" swrid="5117103" athleteid="2064">
              <RESULTS>
                <RESULT eventid="1075" points="554" reactiontime="+58" swimtime="00:00:25.45" resultid="2065" heatid="2970" lane="5" entrytime="00:00:25.48" entrycourse="LCM" />
                <RESULT eventid="1115" points="538" reactiontime="+70" swimtime="00:01:09.93" resultid="2066" heatid="3010" lane="8" entrytime="00:01:10.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="611" reactiontime="+59" swimtime="00:00:55.28" resultid="2067" heatid="3042" lane="5" entrytime="00:00:56.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nikodem" lastname="Ptak" birthdate="2008-03-27" gender="M" nation="POL" license="100315700396" swrid="5311272" athleteid="2052">
              <RESULTS>
                <RESULT eventid="1075" points="191" reactiontime="+77" swimtime="00:00:36.26" resultid="2053" heatid="2963" lane="4" />
                <RESULT eventid="1139" points="199" reactiontime="+67" swimtime="00:01:20.32" resultid="2054" heatid="3036" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="136" swimtime="00:00:50.44" resultid="2055" heatid="3053" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Werwiński" birthdate="2007-06-07" gender="M" nation="POL" license="100315700404" swrid="5298509" athleteid="2048">
              <RESULTS>
                <RESULT eventid="1075" points="357" reactiontime="+71" swimtime="00:00:29.46" resultid="2049" heatid="2967" lane="1" entrytime="00:00:29.91" entrycourse="LCM" />
                <RESULT eventid="1099" points="292" reactiontime="+77" swimtime="00:00:36.16" resultid="2050" heatid="2991" lane="1" entrytime="00:00:37.66" entrycourse="LCM" />
                <RESULT eventid="1139" points="342" reactiontime="+77" swimtime="00:01:07.05" resultid="2051" heatid="3039" lane="8" entrytime="00:01:07.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Filipiak" birthdate="2003-12-13" gender="M" nation="POL" license="100315700247" swrid="5034215" athleteid="2059">
              <RESULTS>
                <RESULT eventid="1075" points="518" reactiontime="+63" swimtime="00:00:26.02" resultid="2060" heatid="2962" lane="0" />
                <RESULT eventid="1083" points="481" reactiontime="+77" swimtime="00:02:40.92" resultid="2061" heatid="2974" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:18.13" />
                    <SPLIT distance="150" swimtime="00:02:00.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="497" reactiontime="+68" swimtime="00:01:11.79" resultid="2062" heatid="3007" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="508" reactiontime="+63" swimtime="00:00:32.52" resultid="2063" heatid="3050" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+88" swimtime="00:01:53.34" resultid="2094" heatid="2948" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                    <SPLIT distance="100" swimtime="00:00:56.36" />
                    <SPLIT distance="150" swimtime="00:01:27.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2081" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="2029" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="2018" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2059" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+74" swimtime="00:02:00.08" resultid="2095" heatid="2947" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.93" />
                    <SPLIT distance="100" swimtime="00:00:56.83" />
                    <SPLIT distance="150" swimtime="00:01:26.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2085" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2068" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="2088" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2022" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="1656" name="KS Warta Poznań">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Szymkowiak" birthdate="1980-04-12" gender="M" nation="POL" license="500115700523" swrid="5312534" athleteid="1748">
              <RESULTS>
                <RESULT eventid="1075" points="501" reactiontime="+76" swimtime="00:00:26.32" resultid="1749" heatid="2962" lane="6" />
                <RESULT eventid="1115" points="601" reactiontime="+68" swimtime="00:01:07.38" resultid="1750" heatid="3006" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="620" reactiontime="+74" swimtime="00:00:30.42" resultid="1751" heatid="3052" lane="4" />
                <RESULT eventid="1171" points="461" reactiontime="+79" swimtime="00:02:27.57" resultid="1752" heatid="3069" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="100" swimtime="00:01:12.64" />
                    <SPLIT distance="150" swimtime="00:01:54.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Kolańczyk" birthdate="2006-09-05" gender="F" nation="POL" license="100115600428" swrid="5162144" athleteid="1666">
              <RESULTS>
                <RESULT eventid="1071" points="601" swimtime="00:00:28.04" resultid="1667" heatid="2959" lane="2" entrytime="00:00:27.71" entrycourse="LCM" />
                <RESULT eventid="1087" points="559" reactiontime="+79" swimtime="00:01:07.33" resultid="1668" heatid="2979" lane="9" entrytime="00:01:08.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="537" reactiontime="+68" swimtime="00:00:30.05" resultid="1669" heatid="3016" lane="6" entrytime="00:00:29.70" entrycourse="LCM" />
                <RESULT eventid="1135" points="599" reactiontime="+69" swimtime="00:01:01.33" resultid="1670" heatid="3034" lane="7" entrytime="00:01:01.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Smektała" birthdate="2004-04-15" gender="F" nation="POL" license="100115600586" swrid="5114691" athleteid="1815">
              <RESULTS>
                <RESULT eventid="1087" points="587" reactiontime="+76" swimtime="00:01:06.26" resultid="1816" heatid="2979" lane="3" entrytime="00:01:06.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="518" swimtime="00:00:30.41" resultid="1817" heatid="3016" lane="2" entrytime="00:00:29.80" entrycourse="LCM" />
                <RESULT eventid="1151" points="542" reactiontime="+70" swimtime="00:02:29.34" resultid="1818" heatid="3058" lane="4" entrytime="00:02:30.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:11.98" />
                    <SPLIT distance="150" swimtime="00:01:50.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Derek" birthdate="2004-01-30" gender="M" nation="POL" license="100115700568" swrid="5034148" athleteid="1770">
              <RESULTS>
                <RESULT eventid="1075" points="419" swimtime="00:00:27.94" resultid="1771" heatid="2968" lane="2" entrytime="00:00:28.12" entrycourse="LCM" />
                <RESULT eventid="1107" points="467" reactiontime="+73" swimtime="00:02:11.40" resultid="1772" heatid="3000" lane="5" entrytime="00:02:12.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="100" swimtime="00:01:03.64" />
                    <SPLIT distance="150" swimtime="00:01:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="489" reactiontime="+71" swimtime="00:00:59.54" resultid="1773" heatid="3040" lane="6" entrytime="00:01:00.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwier" lastname="Cichocki" birthdate="2004-06-04" gender="M" nation="POL" license="100115700247" swrid="5034130" athleteid="1796">
              <RESULTS>
                <RESULT eventid="1083" points="528" reactiontime="+72" swimtime="00:02:36.03" resultid="1797" heatid="2976" lane="5" entrytime="00:02:30.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:18.95" />
                    <SPLIT distance="150" swimtime="00:01:59.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="509" reactiontime="+71" swimtime="00:01:11.22" resultid="1798" heatid="3010" lane="3" entrytime="00:01:08.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="536" reactiontime="+71" swimtime="00:00:31.94" resultid="1799" heatid="3057" lane="7" entrytime="00:00:31.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oleksandr" lastname="Kuchuk" birthdate="1986-06-26" gender="M" nation="POL" license="500115700583" swrid="5435202" athleteid="1781">
              <RESULTS>
                <RESULT eventid="1083" points="438" reactiontime="+78" swimtime="00:02:46.07" resultid="1782" heatid="2975" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:15.89" />
                    <SPLIT distance="150" swimtime="00:02:00.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="492" reactiontime="+75" swimtime="00:01:12.04" resultid="1783" heatid="3007" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="520" reactiontime="+74" swimtime="00:00:32.25" resultid="1784" heatid="3053" lane="4" />
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="1785" heatid="3070" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Zajączek" birthdate="1976-07-17" gender="F" nation="POL" license="500115600524" swrid="5455051" athleteid="1774">
              <RESULTS>
                <RESULT eventid="1079" points="147" swimtime="00:04:23.37" resultid="1775" heatid="2972" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.48" />
                    <SPLIT distance="100" swimtime="00:02:08.02" />
                    <SPLIT distance="150" swimtime="00:03:15.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustaw" lastname="Warzocha" birthdate="2004-09-21" gender="M" nation="POL" license="100115700587" swrid="5034133" athleteid="1804">
              <RESULTS>
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="1805" heatid="2974" lane="5" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="1806" heatid="3043" lane="1" entrytime="00:00:55.19" entrycourse="LCM" />
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="1807" heatid="3072" lane="4" entrytime="00:02:13.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Malwina" lastname="Mikołajczak" birthdate="2006-11-16" gender="F" nation="POL" license="100115600419" swrid="5071600" athleteid="1712">
              <RESULTS>
                <RESULT eventid="1071" points="559" reactiontime="+55" swimtime="00:00:28.72" resultid="1713" heatid="2958" lane="5" entrytime="00:00:28.51" entrycourse="LCM" />
                <RESULT eventid="1095" points="565" reactiontime="+79" swimtime="00:00:32.63" resultid="1714" heatid="2987" lane="7" entrytime="00:00:32.21" entrycourse="LCM" />
                <RESULT eventid="1127" points="565" reactiontime="+75" swimtime="00:02:29.18" resultid="1715" heatid="3026" lane="4" entrytime="00:02:29.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                    <SPLIT distance="150" swimtime="00:01:52.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="587" reactiontime="+73" swimtime="00:01:08.75" resultid="1716" heatid="3062" lane="2" entrytime="00:01:09.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Celmer" birthdate="2003-12-28" gender="F" nation="POL" license="100115600361" swrid="4940377" athleteid="1692">
              <RESULTS>
                <RESULT eventid="1071" points="717" reactiontime="+71" swimtime="00:00:26.44" resultid="1693" heatid="2953" lane="7" />
                <RESULT eventid="1119" points="666" reactiontime="+65" swimtime="00:00:27.97" resultid="1694" heatid="3016" lane="4" entrytime="00:00:27.80" entrycourse="LCM" />
                <RESULT eventid="1135" points="724" reactiontime="+70" swimtime="00:00:57.57" resultid="1695" heatid="3034" lane="4" entrytime="00:00:57.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Baranowska" birthdate="2003-06-13" gender="F" nation="POL" license="100115600359" swrid="4995068" athleteid="1696">
              <RESULTS>
                <RESULT eventid="1071" points="578" reactiontime="+78" swimtime="00:00:28.41" resultid="1697" heatid="2958" lane="3" entrytime="00:00:28.61" entrycourse="LCM" />
                <RESULT eventid="1103" points="573" reactiontime="+74" swimtime="00:02:15.96" resultid="1698" heatid="2997" lane="0" entrytime="00:02:19.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:05.34" />
                    <SPLIT distance="150" swimtime="00:01:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="587" reactiontime="+70" swimtime="00:01:01.73" resultid="1699" heatid="3033" lane="5" entrytime="00:01:02.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Zadorożny" birthdate="1978-08-31" gender="M" nation="POL" license="500115700461" swrid="4920304" athleteid="1768">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="1769" heatid="2961" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olaf" lastname="Kosiorek" birthdate="2007-06-15" gender="M" nation="POL" license="100115700483" swrid="4838389" athleteid="1756">
              <RESULTS>
                <RESULT eventid="1075" points="363" reactiontime="+75" swimtime="00:00:29.30" resultid="1757" heatid="2968" lane="9" entrytime="00:00:29.10" entrycourse="LCM" />
                <RESULT eventid="1139" points="418" reactiontime="+65" swimtime="00:01:02.73" resultid="1758" heatid="3039" lane="5" entrytime="00:01:03.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Wrzeszczyńska" birthdate="2007-07-03" gender="F" nation="POL" license="100115600456" swrid="5162152" athleteid="1676">
              <RESULTS>
                <RESULT eventid="1071" points="598" reactiontime="+78" swimtime="00:00:28.08" resultid="1677" heatid="2959" lane="6" entrytime="00:00:27.62" entrycourse="LCM" />
                <RESULT eventid="1119" points="531" reactiontime="+74" swimtime="00:00:30.16" resultid="1678" heatid="3016" lane="0" entrytime="00:00:30.10" entrycourse="LCM" />
                <RESULT eventid="1159" points="489" reactiontime="+75" swimtime="00:01:13.07" resultid="1679" heatid="3061" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julian" lastname="Januszewski" birthdate="2007-04-16" gender="M" nation="POL" license="100115700478" swrid="4838390" athleteid="1845">
              <RESULTS>
                <RESULT eventid="1099" points="334" reactiontime="+59" swimtime="00:00:34.59" resultid="1846" heatid="2991" lane="5" entrytime="00:00:35.35" entrycourse="LCM" />
                <RESULT eventid="1163" points="322" reactiontime="+74" swimtime="00:01:15.61" resultid="1847" heatid="3064" lane="6" entrytime="00:01:17.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Kotecka" birthdate="1965-05-08" gender="F" nation="POL" license="100115600357" swrid="4754727" athleteid="1852">
              <RESULTS>
                <RESULT eventid="1103" points="208" reactiontime="+101" swimtime="00:03:10.44" resultid="1853" heatid="2995" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                    <SPLIT distance="100" swimtime="00:01:30.99" />
                    <SPLIT distance="150" swimtime="00:02:21.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="180" reactiontime="+137" swimtime="00:03:38.45" resultid="1854" heatid="3025" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.89" />
                    <SPLIT distance="100" swimtime="00:01:48.42" />
                    <SPLIT distance="150" swimtime="00:02:44.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="198" swimtime="00:01:28.68" resultid="1855" heatid="3029" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="217" reactiontime="+103" swimtime="00:06:33.14" resultid="1856" heatid="3073" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                    <SPLIT distance="100" swimtime="00:01:33.46" />
                    <SPLIT distance="150" swimtime="00:02:24.64" />
                    <SPLIT distance="200" swimtime="00:03:15.99" />
                    <SPLIT distance="250" swimtime="00:04:07.21" />
                    <SPLIT distance="300" swimtime="00:04:58.23" />
                    <SPLIT distance="350" swimtime="00:05:47.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Thiem" birthdate="1963-02-17" gender="M" nation="POL" license="100115700345" swrid="4754725" athleteid="1819">
              <RESULTS>
                <RESULT eventid="1091" points="165" swimtime="00:01:30.20" resultid="1820" heatid="2980" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="158" reactiontime="+104" swimtime="00:03:08.38" resultid="1821" heatid="2998" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                    <SPLIT distance="100" swimtime="00:01:32.55" />
                    <SPLIT distance="150" swimtime="00:02:21.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sylwia" lastname="Gorockiewicz" birthdate="1975-03-29" gender="F" nation="POL" license="500115600525" swrid="4837788" athleteid="1685">
              <RESULTS>
                <RESULT eventid="1071" points="68" reactiontime="+109" swimtime="00:00:57.98" resultid="1686" heatid="2953" lane="0" />
                <RESULT eventid="1079" points="110" reactiontime="+116" swimtime="00:04:49.61" resultid="1687" heatid="2972" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.52" />
                    <SPLIT distance="100" swimtime="00:02:18.97" />
                    <SPLIT distance="150" swimtime="00:03:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="98" reactiontime="+104" swimtime="00:02:18.65" resultid="1688" heatid="3003" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Szczepańska" birthdate="2003-09-06" gender="F" nation="POL" license="100115600375" swrid="5030844" athleteid="1857">
              <RESULTS>
                <RESULT eventid="1103" points="649" reactiontime="+80" swimtime="00:02:10.45" resultid="1858" heatid="2997" lane="4" entrytime="00:02:11.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                    <SPLIT distance="100" swimtime="00:01:04.33" />
                    <SPLIT distance="150" swimtime="00:01:38.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="662" reactiontime="+75" swimtime="00:00:59.31" resultid="1859" heatid="3034" lane="5" entrytime="00:00:59.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="652" reactiontime="+80" swimtime="00:04:32.68" resultid="1860" heatid="3074" lane="4" entrytime="00:04:39.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:06.17" />
                    <SPLIT distance="150" swimtime="00:01:41.26" />
                    <SPLIT distance="200" swimtime="00:02:16.15" />
                    <SPLIT distance="250" swimtime="00:02:50.87" />
                    <SPLIT distance="300" swimtime="00:03:25.55" />
                    <SPLIT distance="350" swimtime="00:04:00.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Matysiak" birthdate="2003-02-22" gender="M" nation="POL" license="100115700367" swrid="4940370" athleteid="1848">
              <RESULTS>
                <RESULT eventid="1099" points="506" reactiontime="+57" swimtime="00:00:30.10" resultid="1849" heatid="2993" lane="0" entrytime="00:00:29.32" entrycourse="LCM" />
                <RESULT eventid="1131" status="DNS" swimtime="00:00:00.00" resultid="1850" heatid="3027" lane="5" entrytime="00:02:21.60" entrycourse="LCM" />
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="1851" heatid="3072" lane="2" entrytime="00:02:20.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matylda" lastname="Kaniasta" birthdate="2005-05-16" gender="F" nation="POL" license="100115600541" swrid="4981607" athleteid="1708">
              <RESULTS>
                <RESULT eventid="1071" points="434" reactiontime="+90" swimtime="00:00:31.26" resultid="1709" heatid="2956" lane="9" entrytime="00:00:31.34" entrycourse="LCM" />
                <RESULT eventid="1103" points="440" reactiontime="+82" swimtime="00:02:28.49" resultid="1710" heatid="2996" lane="1" entrytime="00:02:33.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:08.97" />
                    <SPLIT distance="150" swimtime="00:01:48.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="433" reactiontime="+77" swimtime="00:01:08.35" resultid="1711" heatid="3032" lane="0" entrytime="00:01:08.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Kordalska" birthdate="2008-03-24" gender="F" nation="POL" license="100115600503" swrid="4416124" athleteid="1812">
              <RESULTS>
                <RESULT eventid="1087" points="398" reactiontime="+69" swimtime="00:01:15.38" resultid="1813" heatid="2977" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="400" reactiontime="+64" swimtime="00:00:33.13" resultid="1814" heatid="3014" lane="3" entrytime="00:00:34.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kajetan" lastname="Krucki" birthdate="2006-09-16" gender="M" nation="POL" license="100115700431" swrid="5162145" athleteid="1837">
              <RESULTS>
                <RESULT eventid="1099" points="579" reactiontime="+70" swimtime="00:00:28.79" resultid="1838" heatid="2993" lane="8" entrytime="00:00:29.23" entrycourse="LCM" />
                <RESULT eventid="1123" points="584" reactiontime="+67" swimtime="00:00:26.64" resultid="1839" heatid="3024" lane="8" entrytime="00:00:26.49" entrycourse="LCM" />
                <RESULT eventid="1139" points="599" reactiontime="+63" swimtime="00:00:55.63" resultid="1840" heatid="3042" lane="3" entrytime="00:00:56.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Witt" birthdate="1991-08-11" gender="M" nation="POL" license="500115700645" swrid="5062813" athleteid="1720">
              <RESULTS>
                <RESULT eventid="1075" points="544" reactiontime="+76" swimtime="00:00:25.61" resultid="1721" heatid="2964" lane="1" />
                <RESULT eventid="1107" points="438" reactiontime="+76" swimtime="00:02:14.30" resultid="1722" heatid="2998" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:03.29" />
                    <SPLIT distance="150" swimtime="00:01:39.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="499" reactiontime="+76" swimtime="00:00:28.06" resultid="1723" heatid="3018" lane="9" />
                <RESULT eventid="1139" points="557" reactiontime="+76" swimtime="00:00:56.99" resultid="1724" heatid="3036" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Wróbel" birthdate="2007-10-20" gender="M" nation="POL" license="100115700476" swrid="4838417" athleteid="1789">
              <RESULTS>
                <RESULT eventid="1083" points="332" reactiontime="+80" swimtime="00:03:02.08" resultid="1790" heatid="2976" lane="9" entrytime="00:03:06.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:26.29" />
                    <SPLIT distance="150" swimtime="00:02:14.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="316" reactiontime="+73" swimtime="00:00:38.06" resultid="1791" heatid="3055" lane="4" entrytime="00:00:38.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Chybiński" birthdate="2008-09-06" gender="M" nation="POL" license="100115700500" swrid="4997017" athleteid="1753">
              <RESULTS>
                <RESULT eventid="1075" points="435" reactiontime="+83" swimtime="00:00:27.59" resultid="1754" heatid="2968" lane="4" entrytime="00:00:27.55" entrycourse="LCM" />
                <RESULT eventid="1139" points="449" reactiontime="+89" swimtime="00:01:01.24" resultid="1755" heatid="3041" lane="9" entrytime="00:00:59.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Waraczewski" birthdate="1962-04-19" gender="M" nation="POL" license="100115700344" swrid="4992781" athleteid="1786">
              <RESULTS>
                <RESULT eventid="1083" points="245" reactiontime="+93" swimtime="00:03:21.41" resultid="1787" heatid="2974" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                    <SPLIT distance="100" swimtime="00:01:34.98" />
                    <SPLIT distance="150" swimtime="00:02:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="238" reactiontime="+87" swimtime="00:01:31.73" resultid="1788" heatid="3006" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Celmer" birthdate="2007-03-26" gender="F" nation="POL" license="100115600449" swrid="5162156" athleteid="1825">
              <RESULTS>
                <RESULT eventid="1095" points="652" reactiontime="+77" swimtime="00:00:31.11" resultid="1826" heatid="2987" lane="3" entrytime="00:00:31.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Błażej" lastname="Wachowski" birthdate="1980-10-08" gender="M" nation="POL" license="100115700545" swrid="4595659" athleteid="1861">
              <RESULTS>
                <RESULT eventid="1107" points="338" reactiontime="+98" swimtime="00:02:26.41" resultid="1862" heatid="2999" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:09.77" />
                    <SPLIT distance="150" swimtime="00:01:47.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="257" reactiontime="+95" swimtime="00:02:54.10" resultid="1863" heatid="3059" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:18.86" />
                    <SPLIT distance="150" swimtime="00:02:05.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="322" reactiontime="+88" swimtime="00:05:21.00" resultid="1864" heatid="3076" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:15.32" />
                    <SPLIT distance="150" swimtime="00:01:56.64" />
                    <SPLIT distance="200" swimtime="00:02:37.91" />
                    <SPLIT distance="250" swimtime="00:03:19.44" />
                    <SPLIT distance="300" swimtime="00:04:01.12" />
                    <SPLIT distance="350" swimtime="00:04:42.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Budny" birthdate="2006-05-04" gender="M" nation="POL" license="100115700424" swrid="5162174" athleteid="1657">
              <RESULTS>
                <RESULT eventid="1067" points="498" reactiontime="+64" swimtime="00:05:07.56" resultid="1658" heatid="2950" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="100" swimtime="00:01:09.56" />
                    <SPLIT distance="150" swimtime="00:01:49.33" />
                    <SPLIT distance="200" swimtime="00:02:29.34" />
                    <SPLIT distance="250" swimtime="00:03:10.25" />
                    <SPLIT distance="300" swimtime="00:03:54.55" />
                    <SPLIT distance="350" swimtime="00:04:32.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="508" reactiontime="+72" swimtime="00:00:30.07" resultid="1659" heatid="2992" lane="6" entrytime="00:00:29.90" entrycourse="LCM" />
                <RESULT eventid="1147" points="507" reactiontime="+65" swimtime="00:00:32.53" resultid="1660" heatid="3056" lane="5" entrytime="00:00:32.80" entrycourse="LCM" />
                <RESULT eventid="1171" points="492" reactiontime="+65" swimtime="00:02:24.33" resultid="1661" heatid="3072" lane="1" entrytime="00:02:22.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:08.17" />
                    <SPLIT distance="150" swimtime="00:01:50.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Volodymyr" lastname="Kuz" birthdate="2005-03-16" gender="M" nation="POL" license="100115700540" swrid="5198883" athleteid="1800">
              <RESULTS>
                <RESULT eventid="1083" points="459" reactiontime="+81" swimtime="00:02:43.42" resultid="1801" heatid="2976" lane="8" entrytime="00:02:45.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:17.94" />
                    <SPLIT distance="150" swimtime="00:02:01.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="482" reactiontime="+81" swimtime="00:01:12.54" resultid="1802" heatid="3009" lane="6" entrytime="00:01:12.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="495" reactiontime="+73" swimtime="00:00:32.80" resultid="1803" heatid="3057" lane="0" entrytime="00:00:32.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Kuca" birthdate="1994-07-23" gender="M" nation="POL" license="100115700396" swrid="4213120" athleteid="1725">
              <RESULTS>
                <RESULT eventid="1075" points="617" reactiontime="+72" swimtime="00:00:24.55" resultid="1726" heatid="2964" lane="4" />
                <RESULT eventid="1171" points="572" reactiontime="+64" swimtime="00:02:17.33" resultid="1727" heatid="3071" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.25" />
                    <SPLIT distance="100" swimtime="00:01:04.12" />
                    <SPLIT distance="150" swimtime="00:01:45.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Chruściel" birthdate="2007-04-23" gender="M" nation="POL" license="100115700450" swrid="5162166" athleteid="1841">
              <RESULTS>
                <RESULT eventid="1099" points="360" reactiontime="+65" swimtime="00:00:33.72" resultid="1842" heatid="2990" lane="8" />
                <RESULT eventid="1123" points="361" reactiontime="+73" swimtime="00:00:31.25" resultid="1843" heatid="3022" lane="9" entrytime="00:00:31.53" entrycourse="LCM" />
                <RESULT eventid="1147" points="334" reactiontime="+70" swimtime="00:00:37.40" resultid="1844" heatid="3051" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Krasowski" birthdate="2006-10-12" gender="M" nation="POL" license="100115700430" swrid="5162163" athleteid="1876">
              <RESULTS>
                <RESULT eventid="1115" points="503" reactiontime="+69" swimtime="00:01:11.52" resultid="1877" heatid="3009" lane="5" entrytime="00:01:10.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="491" reactiontime="+66" swimtime="00:00:32.88" resultid="1878" heatid="3056" lane="6" entrytime="00:00:33.06" entrycourse="LCM" />
                <RESULT eventid="1171" points="482" reactiontime="+69" swimtime="00:02:25.35" resultid="1879" heatid="3072" lane="8" entrytime="00:02:26.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:11.32" />
                    <SPLIT distance="150" swimtime="00:01:52.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Dopieralski" birthdate="2010-04-18" gender="M" nation="POL" license="100115700628" swrid="5278387" athleteid="1762">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="1763" heatid="2963" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Krupińska" birthdate="1953-05-24" gender="F" nation="POL" license="500115600520" swrid="4992790" athleteid="1680">
              <RESULTS>
                <RESULT eventid="1071" points="107" reactiontime="+111" swimtime="00:00:49.85" resultid="1681" heatid="2953" lane="5" />
                <RESULT eventid="1079" points="155" reactiontime="+107" swimtime="00:04:18.78" resultid="1682" heatid="2972" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.44" />
                    <SPLIT distance="100" swimtime="00:02:06.26" />
                    <SPLIT distance="150" swimtime="00:03:13.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="152" reactiontime="+127" swimtime="00:02:00.01" resultid="1683" heatid="3003" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="169" reactiontime="+90" swimtime="00:00:53.12" resultid="1684" heatid="3044" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Szukała" birthdate="2003-09-23" gender="M" nation="POL" license="100115700376" swrid="5004231" athleteid="1792">
              <RESULTS>
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="1793" heatid="2976" lane="7" entrytime="00:02:41.84" entrycourse="LCM" />
                <RESULT eventid="1115" status="DNS" swimtime="00:00:00.00" resultid="1794" heatid="3009" lane="2" entrytime="00:01:12.74" entrycourse="LCM" />
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="1795" heatid="3057" lane="8" entrytime="00:00:31.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Czechyra" birthdate="2006-08-04" gender="F" nation="POL" license="100115600413" swrid="5135298" athleteid="1704">
              <RESULTS>
                <RESULT eventid="1071" points="409" swimtime="00:00:31.88" resultid="1705" heatid="2956" lane="2" entrytime="00:00:30.77" entrycourse="LCM" />
                <RESULT eventid="1103" points="413" swimtime="00:02:31.66" resultid="1706" heatid="2996" lane="2" entrytime="00:02:31.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:53.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="419" reactiontime="+68" swimtime="00:01:09.07" resultid="1707" heatid="3031" lane="4" entrytime="00:01:09.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Czechyra" birthdate="2003-08-23" gender="F" nation="POL" license="100115600362" swrid="4940375" athleteid="1827">
              <RESULTS>
                <RESULT eventid="1095" points="547" reactiontime="+74" swimtime="00:00:32.98" resultid="1828" heatid="2987" lane="2" entrytime="00:00:32.07" entrycourse="LCM" />
                <RESULT eventid="1103" points="540" reactiontime="+77" swimtime="00:02:18.69" resultid="1829" heatid="2997" lane="5" entrytime="00:02:11.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:08.14" />
                    <SPLIT distance="150" swimtime="00:01:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="545" reactiontime="+75" swimtime="00:02:31.01" resultid="1830" heatid="3025" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:14.95" />
                    <SPLIT distance="150" swimtime="00:01:53.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="584" reactiontime="+77" swimtime="00:01:08.84" resultid="1831" heatid="3062" lane="3" entrytime="00:01:08.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Kuśnierczak" birthdate="2008-01-26" gender="F" nation="POL" license="100115600506" swrid="4998018" athleteid="1873">
              <RESULTS>
                <RESULT eventid="1111" points="417" reactiontime="+83" swimtime="00:01:25.78" resultid="1874" heatid="3004" lane="6" entrytime="00:01:26.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="453" reactiontime="+76" swimtime="00:00:38.26" resultid="1875" heatid="3048" lane="2" entrytime="00:00:39.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Szafrański" birthdate="2007-02-01" gender="M" nation="POL" license="100115700479" swrid="4997918" athleteid="1759">
              <RESULTS>
                <RESULT eventid="1075" points="436" reactiontime="+69" swimtime="00:00:27.57" resultid="1760" heatid="2969" lane="0" entrytime="00:00:27.52" entrycourse="LCM" />
                <RESULT eventid="1147" points="484" reactiontime="+71" swimtime="00:00:33.04" resultid="1761" heatid="3056" lane="3" entrytime="00:00:32.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Rybak" birthdate="2007-04-23" gender="F" nation="POL" license="100115600454" swrid="5162165" athleteid="1671">
              <RESULTS>
                <RESULT eventid="1071" points="565" reactiontime="+61" swimtime="00:00:28.63" resultid="1672" heatid="2952" lane="0" />
                <RESULT eventid="1095" points="548" reactiontime="+62" swimtime="00:00:32.95" resultid="1673" heatid="2984" lane="6" />
                <RESULT eventid="1119" points="520" reactiontime="+55" swimtime="00:00:30.37" resultid="1674" heatid="3015" lane="7" entrytime="00:00:31.53" entrycourse="LCM" />
                <RESULT eventid="1143" points="545" reactiontime="+63" swimtime="00:00:35.99" resultid="1675" heatid="3049" lane="6" entrytime="00:00:35.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Chudy" birthdate="1997-06-21" gender="M" nation="POL" license="100115700495" swrid="4286914" athleteid="1822">
              <RESULTS>
                <RESULT eventid="1091" points="747" reactiontime="+72" swimtime="00:00:54.54" resultid="1823" heatid="2982" lane="4" entrytime="00:00:53.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="729" reactiontime="+74" swimtime="00:00:24.74" resultid="1824" heatid="3024" lane="4" entrytime="00:00:23.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Gryko" birthdate="2009-06-03" gender="F" nation="POL" license="100115600557" swrid="5198903" athleteid="1776">
              <RESULTS>
                <RESULT eventid="1079" points="385" reactiontime="+79" swimtime="00:03:11.11" resultid="1777" heatid="2973" lane="8" entrytime="00:03:07.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:30.85" />
                    <SPLIT distance="150" swimtime="00:02:21.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="385" reactiontime="+70" swimtime="00:01:28.15" resultid="1778" heatid="3004" lane="3" entrytime="00:01:26.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="404" reactiontime="+62" swimtime="00:00:39.76" resultid="1779" heatid="3045" lane="0" />
                <RESULT eventid="1167" points="443" reactiontime="+71" swimtime="00:02:45.32" resultid="1780" heatid="3067" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:19.41" />
                    <SPLIT distance="150" swimtime="00:02:07.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Meyer" birthdate="2005-08-08" gender="M" nation="POL" license="100115700494" swrid="5179173" athleteid="1764">
              <RESULTS>
                <RESULT eventid="1075" points="499" reactiontime="+79" swimtime="00:00:26.35" resultid="1765" heatid="2964" lane="8" />
                <RESULT eventid="1099" points="507" reactiontime="+64" swimtime="00:00:30.08" resultid="1766" heatid="2992" lane="3" entrytime="00:00:29.86" entrycourse="LCM" />
                <RESULT eventid="1163" points="475" reactiontime="+62" swimtime="00:01:06.43" resultid="1767" heatid="3065" lane="1" entrytime="00:01:05.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Ławrynowicz" birthdate="2003-07-31" gender="F" nation="POL" license="100115600569" swrid="4797472" athleteid="1700">
              <RESULTS>
                <RESULT eventid="1071" points="504" reactiontime="+76" swimtime="00:00:29.73" resultid="1701" heatid="2957" lane="4" entrytime="00:00:29.39" entrycourse="LCM" />
                <RESULT eventid="1103" points="516" reactiontime="+78" swimtime="00:02:20.84" resultid="1702" heatid="2995" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:08.06" />
                    <SPLIT distance="150" swimtime="00:01:44.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="506" reactiontime="+68" swimtime="00:01:04.85" resultid="1703" heatid="3033" lane="0" entrytime="00:01:04.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Skolasiński" birthdate="2005-03-09" gender="M" nation="POL" license="100115700391" swrid="5084033" athleteid="1662">
              <RESULTS>
                <RESULT eventid="1067" points="573" reactiontime="+83" swimtime="00:04:53.48" resultid="1663" heatid="2950" lane="4" entrytime="00:04:46.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="100" swimtime="00:01:04.74" />
                    <SPLIT distance="150" swimtime="00:01:44.88" />
                    <SPLIT distance="200" swimtime="00:02:24.81" />
                    <SPLIT distance="250" swimtime="00:03:04.18" />
                    <SPLIT distance="300" swimtime="00:03:44.88" />
                    <SPLIT distance="350" swimtime="00:04:19.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="563" reactiontime="+82" swimtime="00:00:31.41" resultid="1664" heatid="3057" lane="6" entrytime="00:00:30.84" entrycourse="LCM" />
                <RESULT eventid="1171" points="589" reactiontime="+75" swimtime="00:02:15.93" resultid="1665" heatid="3072" lane="5" entrytime="00:02:15.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:01:08.75" />
                    <SPLIT distance="150" swimtime="00:01:45.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Kosiedowski" birthdate="1979-01-02" gender="M" nation="POL" license="500115700566" athleteid="1733">
              <RESULTS>
                <RESULT eventid="1075" points="271" reactiontime="+91" swimtime="00:00:32.28" resultid="1734" heatid="2965" lane="9" />
                <RESULT eventid="1107" points="232" reactiontime="+82" swimtime="00:02:45.83" resultid="1735" heatid="2998" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="150" swimtime="00:02:04.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="243" reactiontime="+76" swimtime="00:00:35.67" resultid="1736" heatid="3017" lane="5" />
                <RESULT eventid="1171" points="213" reactiontime="+78" swimtime="00:03:10.78" resultid="1737" heatid="3069" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:29.53" />
                    <SPLIT distance="150" swimtime="00:02:26.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Janyga" birthdate="1966-03-27" gender="M" nation="POL" license="100115700346" swrid="4992782" athleteid="1832">
              <RESULTS>
                <RESULT eventid="1099" points="379" reactiontime="+75" swimtime="00:00:33.16" resultid="1833" heatid="2990" lane="9" />
                <RESULT eventid="1131" points="295" reactiontime="+87" swimtime="00:02:47.94" resultid="1834" heatid="3028" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="100" swimtime="00:01:23.94" />
                    <SPLIT distance="150" swimtime="00:02:08.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="360" reactiontime="+82" swimtime="00:01:12.86" resultid="1835" heatid="3063" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="302" reactiontime="+94" swimtime="00:05:27.75" resultid="1836" heatid="3075" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:16.44" />
                    <SPLIT distance="150" swimtime="00:01:59.03" />
                    <SPLIT distance="200" swimtime="00:02:42.15" />
                    <SPLIT distance="250" swimtime="00:03:24.93" />
                    <SPLIT distance="300" swimtime="00:04:07.14" />
                    <SPLIT distance="350" swimtime="00:04:48.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Wysocki" birthdate="2004-08-09" gender="M" nation="POL" license="100115700546" swrid="5161574" athleteid="1869">
              <RESULTS>
                <RESULT eventid="1107" points="489" reactiontime="+68" swimtime="00:02:09.44" resultid="1870" heatid="3001" lane="2" entrytime="00:02:06.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                    <SPLIT distance="100" swimtime="00:01:01.58" />
                    <SPLIT distance="150" swimtime="00:01:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="514" reactiontime="+69" swimtime="00:00:58.53" resultid="1871" heatid="3042" lane="7" entrytime="00:00:56.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" status="DNS" swimtime="00:00:00.00" resultid="1872" heatid="3076" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Krzywania" birthdate="2007-04-05" gender="M" nation="POL" license="100115700481" swrid="4838425" athleteid="1880">
              <RESULTS>
                <RESULT eventid="1123" points="408" reactiontime="+73" swimtime="00:00:30.02" resultid="1881" heatid="3022" lane="1" entrytime="00:00:31.39" entrycourse="LCM" />
                <RESULT eventid="1139" points="445" reactiontime="+75" swimtime="00:01:01.44" resultid="1882" heatid="3040" lane="7" entrytime="00:01:02.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antoni" lastname="Bartosik" birthdate="2009-03-12" gender="M" nation="POL" license="100115700563" swrid="5198901" athleteid="1738">
              <RESULTS>
                <RESULT eventid="1075" points="266" reactiontime="+68" swimtime="00:00:32.49" resultid="1739" heatid="2961" lane="0" />
                <RESULT eventid="1115" points="206" reactiontime="+74" swimtime="00:01:36.18" resultid="1740" heatid="3008" lane="8" entrytime="00:01:40.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="210" reactiontime="+73" swimtime="00:00:43.64" resultid="1741" heatid="3051" lane="4" />
                <RESULT eventid="1171" points="260" reactiontime="+68" swimtime="00:02:58.39" resultid="1742" heatid="3071" lane="5" entrytime="00:03:09.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:01:27.66" />
                    <SPLIT distance="150" swimtime="00:02:19.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Ruminiecka" birthdate="2007-08-01" gender="F" nation="POL" license="100115600585" swrid="5002298" athleteid="1689">
              <RESULTS>
                <RESULT eventid="1071" points="472" reactiontime="+72" swimtime="00:00:30.38" resultid="1690" heatid="2956" lane="4" entrytime="00:00:30.16" entrycourse="LCM" />
                <RESULT eventid="1135" points="452" reactiontime="+67" swimtime="00:01:07.33" resultid="1691" heatid="3032" lane="1" entrytime="00:01:07.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Bielewicz" birthdate="2005-11-16" gender="M" nation="POL" license="100115700246" swrid="5084123" athleteid="1808">
              <RESULTS>
                <RESULT eventid="1083" points="470" reactiontime="+87" swimtime="00:02:42.16" resultid="1809" heatid="2976" lane="1" entrytime="00:02:44.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:58.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="449" reactiontime="+86" swimtime="00:01:14.25" resultid="1810" heatid="3009" lane="8" entrytime="00:01:15.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="421" reactiontime="+72" swimtime="00:00:34.61" resultid="1811" heatid="3056" lane="1" entrytime="00:00:34.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Lesiński" birthdate="1944-04-13" gender="M" nation="POL" license="500115700616" swrid="4188190" athleteid="1728">
              <RESULTS>
                <RESULT eventid="1075" points="111" reactiontime="+112" swimtime="00:00:43.50" resultid="1729" heatid="2961" lane="5" />
                <RESULT eventid="1099" points="107" reactiontime="+75" swimtime="00:00:50.51" resultid="1730" heatid="2988" lane="1" />
                <RESULT eventid="1139" points="97" reactiontime="+109" swimtime="00:01:42.00" resultid="1731" heatid="3036" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="86" reactiontime="+79" swimtime="00:01:57.09" resultid="1732" heatid="3063" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Makowski" birthdate="2003-08-15" gender="M" nation="POL" license="100115700547" swrid="5150182" athleteid="1865">
              <RESULTS>
                <RESULT eventid="1107" points="554" reactiontime="+84" swimtime="00:02:04.15" resultid="1866" heatid="3001" lane="3" entrytime="00:02:05.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                    <SPLIT distance="100" swimtime="00:01:01.28" />
                    <SPLIT distance="150" swimtime="00:01:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="569" reactiontime="+79" swimtime="00:00:56.60" resultid="1867" heatid="3042" lane="8" entrytime="00:00:56.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="573" reactiontime="+73" swimtime="00:04:24.94" resultid="1868" heatid="3077" lane="4" entrytime="00:04:26.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:03.95" />
                    <SPLIT distance="150" swimtime="00:01:38.13" />
                    <SPLIT distance="200" swimtime="00:02:12.06" />
                    <SPLIT distance="250" swimtime="00:02:46.21" />
                    <SPLIT distance="300" swimtime="00:03:20.21" />
                    <SPLIT distance="350" swimtime="00:03:53.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Życka" birthdate="2007-06-25" gender="F" nation="POL" license="100115600487" swrid="5154995" athleteid="1717">
              <RESULTS>
                <RESULT eventid="1071" points="431" reactiontime="+74" swimtime="00:00:31.32" resultid="1718" heatid="2956" lane="8" entrytime="00:00:31.31" entrycourse="LCM" />
                <RESULT eventid="1135" points="403" reactiontime="+76" swimtime="00:01:09.97" resultid="1719" heatid="3032" lane="7" entrytime="00:01:07.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Chruściel" birthdate="2009-06-19" gender="M" nation="POL" license="100115700554" swrid="5198876" athleteid="1743">
              <RESULTS>
                <RESULT eventid="1075" points="240" reactiontime="+93" swimtime="00:00:33.62" resultid="1744" heatid="2963" lane="2" />
                <RESULT eventid="1139" points="203" reactiontime="+97" swimtime="00:01:19.72" resultid="1745" heatid="3036" lane="2" />
                <RESULT eventid="1147" points="163" swimtime="00:00:47.49" resultid="1746" heatid="3052" lane="5" />
                <RESULT eventid="1171" points="199" reactiontime="+90" swimtime="00:03:15.16" resultid="1747" heatid="3070" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                    <SPLIT distance="100" swimtime="00:01:33.99" />
                    <SPLIT distance="150" swimtime="00:02:33.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+85" swimtime="00:01:44.80" resultid="1883" heatid="2948" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                    <SPLIT distance="100" swimtime="00:00:53.73" />
                    <SPLIT distance="150" swimtime="00:01:20.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1857" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="1764" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="1692" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="1865" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1183" reactiontime="+65" swimtime="00:01:57.93" resultid="1886" heatid="3079" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="100" swimtime="00:01:01.95" />
                    <SPLIT distance="150" swimtime="00:01:31.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1657" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="1837" number="2" />
                    <RELAYPOSITION athleteid="1666" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="1825" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+67" swimtime="00:01:52.19" resultid="1884" heatid="2948" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:00:57.48" />
                    <SPLIT distance="150" swimtime="00:01:25.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1671" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="1841" number="2" />
                    <RELAYPOSITION athleteid="1666" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="1876" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1183" reactiontime="+58" swimtime="00:02:03.75" resultid="1887" heatid="3078" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:04.95" />
                    <SPLIT distance="150" swimtime="00:01:35.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1671" number="1" reactiontime="+58" />
                    <RELAYPOSITION athleteid="1876" number="2" />
                    <RELAYPOSITION athleteid="1841" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="1676" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+60" swimtime="00:01:43.93" resultid="1885" heatid="2947" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.52" />
                    <SPLIT distance="100" swimtime="00:00:50.52" />
                    <SPLIT distance="150" swimtime="00:01:18.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1837" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="1825" number="2" />
                    <RELAYPOSITION athleteid="1676" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="1657" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00304" nation="POL" region="04" clubid="2413" name="TP Zielona Góra">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Karczewski" birthdate="1974-06-11" gender="M" nation="POL" license="100304700490" swrid="5342868" athleteid="2414">
              <RESULTS>
                <RESULT eventid="1075" points="331" reactiontime="+109" swimtime="00:00:30.21" resultid="2415" heatid="2963" lane="9" />
                <RESULT eventid="1091" points="265" reactiontime="+89" swimtime="00:01:16.98" resultid="2416" heatid="2980" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="386" reactiontime="+86" swimtime="00:00:30.57" resultid="2417" heatid="3019" lane="0" />
                <RESULT eventid="1139" points="355" reactiontime="+86" swimtime="00:01:06.19" resultid="2418" heatid="3037" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="15" clubid="2369" name="SMS Poznań">
          <ATHLETES>
            <ATHLETE firstname="Amelia" lastname="Dziadek" birthdate="2005-05-31" gender="F" nation="POL" license="107414600034" swrid="5036198" athleteid="2370">
              <RESULTS>
                <RESULT eventid="1095" points="553" reactiontime="+75" swimtime="00:00:32.87" resultid="2371" heatid="2987" lane="0" entrytime="00:00:32.77" entrycourse="LCM" />
                <RESULT eventid="1127" points="549" reactiontime="+73" swimtime="00:02:30.59" resultid="2372" heatid="3026" lane="5" entrytime="00:02:34.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:12.28" />
                    <SPLIT distance="150" swimtime="00:01:51.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="560" reactiontime="+74" swimtime="00:01:09.81" resultid="2373" heatid="3062" lane="1" entrytime="00:01:09.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00601" nation="POL" region="01" clubid="2717" name="WKS Śląsk">
          <ATHLETES>
            <ATHLETE firstname="Natalia" lastname="Janiszewska" birthdate="2006-05-13" gender="F" nation="POL" license="100601600542" swrid="5113511" athleteid="2718">
              <RESULTS>
                <RESULT eventid="1071" points="604" reactiontime="+77" swimtime="00:00:28.00" resultid="2719" heatid="2959" lane="3" entrytime="00:00:27.54" entrycourse="LCM" />
                <RESULT eventid="1135" points="626" reactiontime="+77" swimtime="00:01:00.44" resultid="2720" heatid="3034" lane="3" entrytime="00:00:59.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Zaremba" birthdate="2005-09-29" gender="M" nation="POL" license="100601700414" swrid="5030685" athleteid="2802">
              <RESULTS>
                <RESULT eventid="1139" points="610" reactiontime="+68" swimtime="00:00:55.31" resultid="2803" heatid="3043" lane="9" entrytime="00:00:55.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="583" reactiontime="+66" swimtime="00:02:16.44" resultid="2804" heatid="3072" lane="3" entrytime="00:02:15.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                    <SPLIT distance="100" swimtime="00:01:07.49" />
                    <SPLIT distance="150" swimtime="00:01:46.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Cebula" birthdate="2003-04-21" gender="M" nation="POL" license="100601700462" swrid="4012910" athleteid="2780">
              <RESULTS>
                <RESULT eventid="1099" points="540" reactiontime="+57" swimtime="00:00:29.46" resultid="2781" heatid="2989" lane="0" />
                <RESULT eventid="1115" points="578" reactiontime="+64" swimtime="00:01:08.27" resultid="2782" heatid="3010" lane="2" entrytime="00:01:09.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="623" reactiontime="+69" swimtime="00:00:30.37" resultid="2783" heatid="3057" lane="3" entrytime="00:00:30.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Dutkowiak" birthdate="2003-10-13" gender="F" nation="POL" license="100601600378" swrid="5023598" athleteid="2721">
              <RESULTS>
                <RESULT eventid="1071" points="555" reactiontime="+81" swimtime="00:00:28.80" resultid="2722" heatid="2958" lane="7" entrytime="00:00:28.82" entrycourse="LCM" />
                <RESULT eventid="1103" points="595" reactiontime="+74" swimtime="00:02:14.29" resultid="2723" heatid="2997" lane="6" entrytime="00:02:14.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:04.60" />
                    <SPLIT distance="150" swimtime="00:01:39.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Szwedzki" birthdate="1994-04-18" gender="M" nation="POL" license="100601700371" swrid="4181303" athleteid="2727">
              <RESULTS>
                <RESULT eventid="1075" points="623" reactiontime="+70" swimtime="00:00:24.47" resultid="2728" heatid="2962" lane="5" />
                <RESULT eventid="1099" points="649" reactiontime="+61" swimtime="00:00:27.72" resultid="2729" heatid="2990" lane="2" />
                <RESULT eventid="1163" points="688" reactiontime="+66" swimtime="00:00:58.72" resultid="2730" heatid="3063" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Głowiak" birthdate="2005-09-20" gender="M" nation="POL" license="100601700429" swrid="5198175" athleteid="2750">
              <RESULTS>
                <RESULT eventid="1083" points="522" reactiontime="+74" swimtime="00:02:36.57" resultid="2751" heatid="2976" lane="6" entrytime="00:02:33.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:16.80" />
                    <SPLIT distance="150" swimtime="00:01:57.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="536" reactiontime="+68" swimtime="00:01:10.01" resultid="2752" heatid="3010" lane="0" entrytime="00:01:10.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="566" swimtime="00:00:31.36" resultid="2753" heatid="3057" lane="2" entrytime="00:00:31.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Bieroński" birthdate="1999-03-23" gender="M" nation="POL" license="100601700350" swrid="4639547" athleteid="2773">
              <RESULTS>
                <RESULT eventid="1099" points="674" reactiontime="+65" swimtime="00:00:27.36" resultid="2774" heatid="2993" lane="5" entrytime="00:00:27.29" entrycourse="LCM" />
                <RESULT eventid="1123" points="627" reactiontime="+79" swimtime="00:00:26.01" resultid="2775" heatid="3024" lane="7" entrytime="00:00:25.95" entrycourse="LCM" />
                <RESULT eventid="1147" points="434" reactiontime="+73" swimtime="00:00:34.25" resultid="2776" heatid="3053" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Pityński" birthdate="2003-09-22" gender="M" nation="POL" license="100601700459" swrid="4979899" athleteid="2793">
              <RESULTS>
                <RESULT eventid="1115" points="593" reactiontime="+66" swimtime="00:01:07.67" resultid="2794" heatid="3010" lane="7" entrytime="00:01:09.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="606" reactiontime="+71" swimtime="00:01:01.24" resultid="2795" heatid="3065" lane="4" entrytime="00:01:01.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Majchrzak" birthdate="2005-03-29" gender="F" nation="POL" license="100601600591" swrid="5166045" athleteid="2760">
              <RESULTS>
                <RESULT eventid="1087" points="571" reactiontime="+80" swimtime="00:01:06.86" resultid="2761" heatid="2979" lane="6" entrytime="00:01:06.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="516" reactiontime="+83" swimtime="00:00:30.44" resultid="2762" heatid="3016" lane="9" entrytime="00:00:30.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Modlińska" birthdate="2005-06-30" gender="F" nation="POL" license="100601600650" swrid="5147673" athleteid="2724">
              <RESULTS>
                <RESULT eventid="1071" points="538" reactiontime="+74" swimtime="00:00:29.09" resultid="2725" heatid="2958" lane="8" entrytime="00:00:28.90" entrycourse="LCM" />
                <RESULT eventid="1103" points="558" reactiontime="+68" swimtime="00:02:17.17" resultid="2726" heatid="2996" lane="5" entrytime="00:02:21.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="100" swimtime="00:01:05.93" />
                    <SPLIT distance="150" swimtime="00:01:42.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Gancarz" birthdate="2003-05-06" gender="F" nation="POL" license="100601600649" swrid="4878929" athleteid="2757">
              <RESULTS>
                <RESULT eventid="1087" points="563" reactiontime="+72" swimtime="00:01:07.18" resultid="2758" heatid="2979" lane="5" entrytime="00:01:06.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="617" reactiontime="+80" swimtime="00:02:12.67" resultid="2759" heatid="2997" lane="3" entrytime="00:02:13.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                    <SPLIT distance="100" swimtime="00:01:04.76" />
                    <SPLIT distance="150" swimtime="00:01:39.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Lipiec" birthdate="2006-04-14" gender="M" nation="POL" license="100601700646" swrid="5166059" athleteid="2744">
              <RESULTS>
                <RESULT eventid="1075" points="566" reactiontime="+65" swimtime="00:00:25.27" resultid="2745" heatid="2971" lane="1" entrytime="00:00:24.94" entrycourse="LCM" />
                <RESULT eventid="1139" points="561" reactiontime="+69" swimtime="00:00:56.86" resultid="2746" heatid="3042" lane="1" entrytime="00:00:56.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kiszczak" birthdate="2000-04-23" gender="M" nation="POL" license="100601700467" swrid="4705231" athleteid="2731">
              <RESULTS>
                <RESULT eventid="1075" points="602" reactiontime="+78" swimtime="00:00:24.76" resultid="2732" heatid="2971" lane="4" entrytime="00:00:23.87" entrycourse="LCM" />
                <RESULT eventid="1099" points="722" reactiontime="+66" swimtime="00:00:26.75" resultid="2733" heatid="2993" lane="4" entrytime="00:00:26.97" entrycourse="LCM" />
                <RESULT eventid="1123" points="672" reactiontime="+73" swimtime="00:00:25.42" resultid="2734" heatid="3024" lane="5" entrytime="00:00:25.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Zawadzka" birthdate="2005-05-28" gender="F" nation="POL" license="100601600448" swrid="5198192" athleteid="2763">
              <RESULTS>
                <RESULT eventid="1087" points="463" reactiontime="+84" swimtime="00:01:11.68" resultid="2764" heatid="2979" lane="7" entrytime="00:01:07.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="555" reactiontime="+72" swimtime="00:00:32.83" resultid="2765" heatid="2987" lane="1" entrytime="00:00:32.23" entrycourse="LCM" />
                <RESULT eventid="1119" points="532" reactiontime="+60" swimtime="00:00:30.14" resultid="2766" heatid="3016" lane="1" entrytime="00:00:30.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Skliński" birthdate="2004-06-14" gender="M" nation="POL" license="100601700411" swrid="5088686" athleteid="2777">
              <RESULTS>
                <RESULT eventid="1099" points="578" reactiontime="+67" swimtime="00:00:28.81" resultid="2778" heatid="2993" lane="2" entrytime="00:00:29.06" entrycourse="LCM" />
                <RESULT eventid="1163" points="543" reactiontime="+70" swimtime="00:01:03.54" resultid="2779" heatid="3065" lane="3" entrytime="00:01:03.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tamara" lastname="Jach" birthdate="2006-09-21" gender="F" nation="POL" license="100601600644" swrid="5166047" athleteid="2784">
              <RESULTS>
                <RESULT eventid="1103" points="585" reactiontime="+69" swimtime="00:02:15.08" resultid="2785" heatid="2995" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:06.27" />
                    <SPLIT distance="150" swimtime="00:01:41.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="548" reactiontime="+80" swimtime="00:00:35.92" resultid="2786" heatid="3049" lane="3" entrytime="00:00:35.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Chyra" birthdate="2003-02-12" gender="F" nation="POL" license="100601600615" swrid="4973970" athleteid="2787">
              <RESULTS>
                <RESULT eventid="1103" points="580" reactiontime="+74" swimtime="00:02:15.44" resultid="2788" heatid="2995" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:41.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="583" reactiontime="+67" swimtime="00:01:08.88" resultid="2789" heatid="3062" lane="6" entrytime="00:01:08.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Rusin" birthdate="2005-01-25" gender="M" nation="POL" license="100601700408" swrid="5088684" athleteid="2799">
              <RESULTS>
                <RESULT eventid="1115" points="425" reactiontime="+80" swimtime="00:01:15.65" resultid="2800" heatid="3009" lane="7" entrytime="00:01:13.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="527" reactiontime="+76" swimtime="00:00:32.12" resultid="2801" heatid="3053" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Klara" lastname="Pityńska" birthdate="2006-02-09" gender="F" nation="POL" license="100601600593" swrid="4995344" athleteid="2754">
              <RESULTS>
                <RESULT eventid="1087" points="461" reactiontime="+84" swimtime="00:01:11.81" resultid="2755" heatid="2978" lane="7" entrytime="00:01:13.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="525" reactiontime="+87" swimtime="00:01:11.32" resultid="2756" heatid="3062" lane="9" entrytime="00:01:11.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cezary" lastname="Leiman" birthdate="2003-03-01" gender="M" nation="POL" license="100601700461" swrid="4979911" athleteid="2735">
              <RESULTS>
                <RESULT eventid="1075" points="515" swimtime="00:00:26.08" resultid="2736" heatid="2970" lane="2" entrytime="00:00:25.64" entrycourse="LCM" />
                <RESULT eventid="1123" points="513" reactiontime="+63" swimtime="00:00:27.81" resultid="2737" heatid="3023" lane="4" entrytime="00:00:27.41" entrycourse="LCM" />
                <RESULT eventid="1139" points="526" reactiontime="+72" swimtime="00:00:58.08" resultid="2738" heatid="3042" lane="4" entrytime="00:00:55.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Hellak" birthdate="2003-03-15" gender="F" nation="POL" license="100601600379" swrid="5023594" athleteid="2747">
              <RESULTS>
                <RESULT eventid="1079" points="599" reactiontime="+80" swimtime="00:02:45.01" resultid="2748" heatid="2973" lane="4" entrytime="00:02:42.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:19.92" />
                    <SPLIT distance="150" swimtime="00:02:02.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="633" swimtime="00:01:00.20" resultid="2749" heatid="3034" lane="2" entrytime="00:01:00.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Stachurski" birthdate="2004-02-27" gender="M" nation="POL" license="100601700590" swrid="4979950" athleteid="2767">
              <RESULTS>
                <RESULT eventid="1091" points="567" reactiontime="+79" swimtime="00:00:59.78" resultid="2768" heatid="2982" lane="2" entrytime="00:01:00.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="607" reactiontime="+59" swimtime="00:04:19.80" resultid="2769" heatid="3077" lane="5" entrytime="00:04:28.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                    <SPLIT distance="100" swimtime="00:01:01.71" />
                    <SPLIT distance="150" swimtime="00:01:34.41" />
                    <SPLIT distance="200" swimtime="00:02:07.61" />
                    <SPLIT distance="250" swimtime="00:02:40.74" />
                    <SPLIT distance="300" swimtime="00:03:14.33" />
                    <SPLIT distance="350" swimtime="00:03:47.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Staszak" birthdate="2004-12-02" gender="M" nation="POL" license="100601700551" swrid="4858850" athleteid="2796">
              <RESULTS>
                <RESULT eventid="1115" points="598" reactiontime="+64" swimtime="00:01:07.48" resultid="2797" heatid="3010" lane="5" entrytime="00:01:08.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="618" reactiontime="+66" swimtime="00:00:26.14" resultid="2798" heatid="3020" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Adamczyk" birthdate="2003-06-02" gender="M" nation="POL" license="100601700376" swrid="5023601" athleteid="2739">
              <RESULTS>
                <RESULT eventid="1075" points="516" reactiontime="+62" swimtime="00:00:26.06" resultid="2740" heatid="2970" lane="1" entrytime="00:00:26.14" entrycourse="LCM" />
                <RESULT eventid="1099" points="526" reactiontime="+57" swimtime="00:00:29.73" resultid="2741" heatid="2993" lane="9" entrytime="00:00:29.52" entrycourse="LCM" />
                <RESULT eventid="1139" points="552" reactiontime="+61" swimtime="00:00:57.18" resultid="2742" heatid="3041" lane="4" entrytime="00:00:57.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="512" reactiontime="+52" swimtime="00:01:04.81" resultid="2743" heatid="3065" lane="2" entrytime="00:01:04.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Lechowska" birthdate="2006-06-13" gender="F" nation="POL" license="100601600643" swrid="5165983" athleteid="2790">
              <RESULTS>
                <RESULT eventid="1111" points="625" reactiontime="+70" swimtime="00:01:14.98" resultid="2791" heatid="3005" lane="4" entrytime="00:01:13.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="581" reactiontime="+69" swimtime="00:02:31.14" resultid="2792" heatid="3068" lane="6" entrytime="00:02:37.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="100" swimtime="00:01:11.17" />
                    <SPLIT distance="150" swimtime="00:01:55.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02202" nation="POL" region="02" clubid="2137" name="MKS ,,Astoria&apos;&apos; Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-13" gender="M" nation="POL" license="102202700126" athleteid="2138">
              <RESULTS>
                <RESULT eventid="1075" points="124" reactiontime="+97" swimtime="00:00:41.84" resultid="2139" heatid="2961" lane="4" />
                <RESULT eventid="1147" points="118" reactiontime="+111" swimtime="00:00:52.86" resultid="2140" heatid="3054" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01016" nation="POL" region="16" clubid="2096" name="MKP Kołobrzeg">
          <ATHLETES>
            <ATHLETE firstname="Natalia" lastname="Szpakiewicz" birthdate="2008-06-29" gender="F" nation="POL" license="101016600085" swrid="5321033" athleteid="2105">
              <RESULTS>
                <RESULT eventid="1071" points="442" reactiontime="+63" swimtime="00:00:31.06" resultid="2106" heatid="2952" lane="6" />
                <RESULT eventid="1119" points="361" reactiontime="+61" swimtime="00:00:34.29" resultid="2107" heatid="3012" lane="1" />
                <RESULT eventid="1135" points="432" reactiontime="+60" swimtime="00:01:08.38" resultid="2108" heatid="3032" lane="8" entrytime="00:01:07.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Głuch" birthdate="2008-06-14" gender="F" nation="POL" license="101016600084" swrid="5321048" athleteid="2097">
              <RESULTS>
                <RESULT eventid="1071" points="455" reactiontime="+78" swimtime="00:00:30.76" resultid="2098" heatid="2955" lane="1" entrytime="00:00:33.14" entrycourse="LCM" />
                <RESULT eventid="1127" points="342" reactiontime="+71" swimtime="00:02:56.24" resultid="2099" heatid="3026" lane="1" entrytime="00:03:05.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="423" swimtime="00:01:08.87" resultid="2100" heatid="3032" lane="2" entrytime="00:01:07.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Jaszewska" birthdate="2008-01-16" gender="F" nation="POL" license="101016600093" swrid="5010042" athleteid="2109">
              <RESULTS>
                <RESULT eventid="1071" points="340" reactiontime="+83" swimtime="00:00:33.89" resultid="2110" heatid="2954" lane="7" entrytime="00:00:36.33" entrycourse="LCM" />
                <RESULT eventid="1135" points="333" reactiontime="+79" swimtime="00:01:14.55" resultid="2111" heatid="3030" lane="4" entrytime="00:01:19.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="280" reactiontime="+62" swimtime="00:00:44.89" resultid="2112" heatid="3047" lane="5" entrytime="00:00:44.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Fedasz" birthdate="2008-01-16" gender="M" nation="POL" license="101016700077" swrid="4790800" athleteid="2117">
              <RESULTS>
                <RESULT eventid="1075" points="403" reactiontime="+69" swimtime="00:00:28.30" resultid="2118" heatid="2967" lane="3" entrytime="00:00:29.56" entrycourse="LCM" />
                <RESULT eventid="1139" points="412" reactiontime="+78" swimtime="00:01:03.03" resultid="2119" heatid="3040" lane="8" entrytime="00:01:02.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="423" reactiontime="+76" swimtime="00:04:53.05" resultid="2120" heatid="3077" lane="2" entrytime="00:04:50.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:09.86" />
                    <SPLIT distance="150" swimtime="00:01:47.43" />
                    <SPLIT distance="200" swimtime="00:02:25.15" />
                    <SPLIT distance="250" swimtime="00:03:02.87" />
                    <SPLIT distance="300" swimtime="00:03:41.95" />
                    <SPLIT distance="350" swimtime="00:04:18.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sara" lastname="Hofman" birthdate="2008-07-29" gender="F" nation="POL" license="101016600094" swrid="4940938" athleteid="2113">
              <RESULTS>
                <RESULT eventid="1071" points="349" reactiontime="+70" swimtime="00:00:33.60" resultid="2114" heatid="2954" lane="5" entrytime="00:00:34.51" entrycourse="LCM" />
                <RESULT eventid="1095" points="301" reactiontime="+77" swimtime="00:00:40.23" resultid="2115" heatid="2986" lane="8" entrytime="00:00:39.10" entrycourse="LCM" />
                <RESULT eventid="1135" points="307" reactiontime="+62" swimtime="00:01:16.57" resultid="2116" heatid="3030" lane="5" entrytime="00:01:19.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Dudała" birthdate="2008-09-06" gender="F" nation="POL" license="101016600103" swrid="5441132" athleteid="2101">
              <RESULTS>
                <RESULT eventid="1071" points="342" reactiontime="+88" swimtime="00:00:33.83" resultid="2102" heatid="2954" lane="3" entrytime="00:00:35.76" entrycourse="LCM" />
                <RESULT eventid="1095" points="273" reactiontime="+76" swimtime="00:00:41.58" resultid="2103" heatid="2986" lane="0" entrytime="00:00:39.97" entrycourse="LCM" />
                <RESULT eventid="1135" points="293" reactiontime="+97" swimtime="00:01:17.83" resultid="2104" heatid="3031" lane="9" entrytime="00:01:17.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00515" nation="POL" region="15" clubid="1442" name="KS Posnania Poznań">
          <ATHLETES>
            <ATHLETE firstname="Zuzanna" lastname="Czech" birthdate="2008-05-29" gender="F" nation="POL" license="100515600290" swrid="5255309" athleteid="1471">
              <RESULTS>
                <RESULT eventid="1071" points="316" reactiontime="+94" swimtime="00:00:34.72" resultid="1472" heatid="2954" lane="4" entrytime="00:00:33.96" entrycourse="LCM" />
                <RESULT eventid="1119" points="225" reactiontime="+90" swimtime="00:00:40.16" resultid="1473" heatid="3014" lane="1" entrytime="00:00:37.63" entrycourse="LCM" />
                <RESULT eventid="1135" points="315" swimtime="00:01:15.96" resultid="1474" heatid="3031" lane="2" entrytime="00:01:15.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Kaczmarek" birthdate="2006-04-17" gender="M" nation="POL" license="100515700239" swrid="5227565" athleteid="1547">
              <RESULTS>
                <RESULT eventid="1083" points="391" reactiontime="+77" swimtime="00:02:52.45" resultid="1548" heatid="2975" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:20.46" />
                    <SPLIT distance="150" swimtime="00:02:06.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="426" reactiontime="+69" swimtime="00:02:15.46" resultid="1549" heatid="3001" lane="0" entrytime="00:02:10.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                    <SPLIT distance="100" swimtime="00:01:03.71" />
                    <SPLIT distance="150" swimtime="00:01:39.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="498" reactiontime="+66" swimtime="00:00:59.15" resultid="1550" heatid="3041" lane="1" entrytime="00:00:59.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Włoch" birthdate="2003-12-02" gender="M" nation="POL" license="100515700178" swrid="5185414" athleteid="1487">
              <RESULTS>
                <RESULT eventid="1075" points="563" reactiontime="+67" swimtime="00:00:25.32" resultid="1488" heatid="2971" lane="7" entrytime="00:00:24.80" entrycourse="LCM" />
                <RESULT eventid="1099" points="404" reactiontime="+66" swimtime="00:00:32.46" resultid="1489" heatid="2989" lane="7" />
                <RESULT eventid="1123" points="494" reactiontime="+63" swimtime="00:00:28.17" resultid="1490" heatid="3024" lane="0" entrytime="00:00:26.86" entrycourse="LCM" />
                <RESULT eventid="1139" points="551" reactiontime="+62" swimtime="00:00:57.20" resultid="1491" heatid="3043" lane="5" entrytime="00:00:54.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Stempak" birthdate="2007-09-08" gender="F" nation="POL" license="100515600269" swrid="5214785" athleteid="1542">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="1543" heatid="2973" lane="0" entrytime="00:03:18.00" entrycourse="LCM" />
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="1544" heatid="3004" lane="7" entrytime="00:01:30.05" entrycourse="LCM" />
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="1545" heatid="3048" lane="1" entrytime="00:00:39.75" entrycourse="LCM" />
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="1546" heatid="3068" lane="8" entrytime="00:03:01.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Kryściak" birthdate="2008-04-01" gender="M" nation="POL" license="100515700286" swrid="5198910" athleteid="1579">
              <RESULTS>
                <RESULT eventid="1091" points="223" reactiontime="+47" swimtime="00:01:21.58" resultid="1580" heatid="2981" lane="1" entrytime="00:01:20.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="240" reactiontime="+55" swimtime="00:00:38.57" resultid="1581" heatid="2989" lane="1" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1123" status="DSQ" swimtime="00:00:00.00" resultid="1582" heatid="3021" lane="7" entrytime="00:00:33.54" entrycourse="LCM" />
                <RESULT eventid="1163" points="235" reactiontime="+56" swimtime="00:01:24.01" resultid="1583" heatid="3064" lane="7" entrytime="00:01:20.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Wielgus" birthdate="2001-03-29" gender="M" nation="POL" license="100515700203" swrid="4905538" athleteid="1505">
              <RESULTS>
                <RESULT eventid="1075" points="510" reactiontime="+69" swimtime="00:00:26.16" resultid="1506" heatid="2970" lane="8" entrytime="00:00:26.25" entrycourse="LCM" />
                <RESULT eventid="1099" points="556" reactiontime="+58" swimtime="00:00:29.17" resultid="1507" heatid="2992" lane="4" entrytime="00:00:29.61" entrycourse="LCM" />
                <RESULT eventid="1163" points="528" reactiontime="+61" swimtime="00:01:04.14" resultid="1508" heatid="3064" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Ćwiertnia" birthdate="2007-08-04" gender="F" nation="POL" license="100515600304" swrid="5198924" athleteid="1475">
              <RESULTS>
                <RESULT eventid="1071" points="385" reactiontime="+59" swimtime="00:00:32.52" resultid="1476" heatid="2955" lane="5" entrytime="00:00:31.88" entrycourse="LCM" />
                <RESULT eventid="1095" points="369" reactiontime="+73" swimtime="00:00:37.60" resultid="1477" heatid="2986" lane="7" entrytime="00:00:37.20" entrycourse="LCM" />
                <RESULT eventid="1127" points="284" reactiontime="+72" swimtime="00:03:07.62" resultid="1478" heatid="3026" lane="7" entrytime="00:02:56.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.60" />
                    <SPLIT distance="150" swimtime="00:02:20.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="295" reactiontime="+68" swimtime="00:01:26.40" resultid="1479" heatid="3061" lane="6" entrytime="00:01:21.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Tomczak" birthdate="2005-01-31" gender="M" nation="POL" license="100515700261" swrid="5384568" athleteid="1497">
              <RESULTS>
                <RESULT eventid="1075" points="432" reactiontime="+70" swimtime="00:00:27.65" resultid="1498" heatid="2968" lane="3" entrytime="00:00:27.65" entrycourse="LCM" />
                <RESULT eventid="1139" points="384" reactiontime="+67" swimtime="00:01:04.49" resultid="1499" heatid="3040" lane="0" entrytime="00:01:02.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Krupiński" birthdate="2003-06-16" gender="M" nation="POL" license="100515700157" swrid="4947332" athleteid="1492">
              <RESULTS>
                <RESULT eventid="1075" points="466" reactiontime="+78" swimtime="00:00:26.97" resultid="1493" heatid="2969" lane="4" entrytime="00:00:26.57" entrycourse="LCM" />
                <RESULT eventid="1107" points="489" reactiontime="+78" swimtime="00:02:09.44" resultid="1494" heatid="3001" lane="7" entrytime="00:02:09.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                    <SPLIT distance="100" swimtime="00:01:02.33" />
                    <SPLIT distance="150" swimtime="00:01:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="525" reactiontime="+79" swimtime="00:00:58.12" resultid="1495" heatid="3041" lane="3" entrytime="00:00:57.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="484" reactiontime="+86" swimtime="00:04:40.28" resultid="1496" heatid="3077" lane="6" entrytime="00:04:42.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:04.87" />
                    <SPLIT distance="150" swimtime="00:01:40.42" />
                    <SPLIT distance="200" swimtime="00:02:16.49" />
                    <SPLIT distance="250" swimtime="00:02:52.72" />
                    <SPLIT distance="300" swimtime="00:03:29.24" />
                    <SPLIT distance="350" swimtime="00:04:05.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Dąbek" birthdate="2005-03-11" gender="F" nation="POL" license="100515600281" swrid="5443305" athleteid="1451">
              <RESULTS>
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="1452" heatid="2956" lane="0" entrytime="00:00:31.33" entrycourse="LCM" />
                <RESULT eventid="1087" points="416" reactiontime="+67" swimtime="00:01:14.27" resultid="1453" heatid="2978" lane="1" entrytime="00:01:13.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="409" reactiontime="+64" swimtime="00:00:32.89" resultid="1454" heatid="3015" lane="8" entrytime="00:00:32.65" entrycourse="LCM" />
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="1455" heatid="3068" lane="1" entrytime="00:02:48.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Zalewski" birthdate="2006-12-06" gender="M" nation="POL" license="100515700253" swrid="4027612" athleteid="1589">
              <RESULTS>
                <RESULT eventid="1107" points="527" reactiontime="+69" swimtime="00:02:06.22" resultid="1590" heatid="2999" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="150" swimtime="00:01:34.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="467" reactiontime="+66" swimtime="00:02:24.20" resultid="1591" heatid="3028" lane="6" entrytime="00:02:26.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:10.00" />
                    <SPLIT distance="150" swimtime="00:01:47.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="512" reactiontime="+66" swimtime="00:00:58.62" resultid="1592" heatid="3036" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Jasnoch" birthdate="2007-10-23" gender="M" nation="POL" license="100515700272" swrid="5198914" athleteid="1584">
              <RESULTS>
                <RESULT eventid="1099" points="303" reactiontime="+78" swimtime="00:00:35.70" resultid="1585" heatid="2991" lane="2" entrytime="00:00:36.04" entrycourse="LCM" />
                <RESULT eventid="1131" points="298" reactiontime="+76" swimtime="00:02:47.40" resultid="1586" heatid="3028" lane="1" entrytime="00:02:44.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:01:20.69" />
                    <SPLIT distance="150" swimtime="00:02:06.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="221" reactiontime="+86" swimtime="00:00:42.92" resultid="1587" heatid="3052" lane="3" />
                <RESULT eventid="1163" points="271" reactiontime="+88" swimtime="00:01:20.04" resultid="1588" heatid="3064" lane="3" entrytime="00:01:16.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Denis" lastname="Osiewicz" birthdate="2008-02-11" gender="M" nation="POL" license="100515700283" swrid="5198906" athleteid="1537">
              <RESULTS>
                <RESULT eventid="1075" points="308" reactiontime="+88" swimtime="00:00:30.96" resultid="1538" heatid="2966" lane="5" entrytime="00:00:30.92" entrycourse="LCM" />
                <RESULT eventid="1091" points="171" reactiontime="+81" swimtime="00:01:29.08" resultid="1539" heatid="2981" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="273" reactiontime="+84" swimtime="00:00:34.32" resultid="1540" heatid="3021" lane="1" entrytime="00:00:33.94" entrycourse="LCM" />
                <RESULT eventid="1139" points="305" reactiontime="+83" swimtime="00:01:09.65" resultid="1541" heatid="3037" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Jagodzińska" birthdate="2008-01-20" gender="F" nation="POL" license="100515600282" swrid="5255316" athleteid="1566">
              <RESULTS>
                <RESULT eventid="1087" points="349" reactiontime="+75" swimtime="00:01:18.79" resultid="1567" heatid="2977" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="380" reactiontime="+70" swimtime="00:00:33.70" resultid="1568" heatid="3014" lane="5" entrytime="00:00:33.91" entrycourse="LCM" />
                <RESULT eventid="1135" points="358" reactiontime="+83" swimtime="00:01:12.77" resultid="1569" heatid="3031" lane="6" entrytime="00:01:13.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olga" lastname="Zarzeczna" birthdate="2005-10-01" gender="F" nation="POL" license="100515600224" swrid="5117085" athleteid="1467">
              <RESULTS>
                <RESULT eventid="1071" points="398" reactiontime="+74" swimtime="00:00:32.17" resultid="1468" heatid="2955" lane="4" entrytime="00:00:31.72" entrycourse="LCM" />
                <RESULT eventid="1103" points="428" reactiontime="+80" swimtime="00:02:29.87" resultid="1469" heatid="2995" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:11.13" />
                    <SPLIT distance="150" swimtime="00:01:51.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="373" reactiontime="+75" swimtime="00:00:40.81" resultid="1470" heatid="3046" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Klimczak" birthdate="2007-10-02" gender="M" nation="POL" license="100515700265" swrid="5198900" athleteid="1518">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="1519" heatid="2961" lane="2" />
                <RESULT eventid="1115" status="DNS" swimtime="00:00:00.00" resultid="1520" heatid="3008" lane="0" />
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="1521" heatid="3052" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Wnuk" birthdate="2001-10-29" gender="M" nation="POL" license="100515700150" swrid="4749884" athleteid="1575">
              <RESULTS>
                <RESULT eventid="1091" points="573" reactiontime="+70" swimtime="00:00:59.57" resultid="1576" heatid="2982" lane="3" entrytime="00:00:59.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="563" reactiontime="+69" swimtime="00:00:26.97" resultid="1577" heatid="3017" lane="6" />
                <RESULT eventid="1155" points="500" reactiontime="+67" swimtime="00:02:19.42" resultid="1578" heatid="3059" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:01:07.01" />
                    <SPLIT distance="150" swimtime="00:01:43.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Bocheńska" birthdate="2005-07-22" gender="F" nation="POL" license="100515600255" swrid="5153525" athleteid="1460">
              <RESULTS>
                <RESULT eventid="1071" points="464" reactiontime="+67" swimtime="00:00:30.57" resultid="1461" heatid="2957" lane="7" entrytime="00:00:29.81" entrycourse="LCM" />
                <RESULT eventid="1135" points="432" reactiontime="+76" swimtime="00:01:08.37" resultid="1462" heatid="3032" lane="3" entrytime="00:01:06.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Nowak" birthdate="2007-02-06" gender="F" nation="POL" license="100515600262" swrid="5087077" athleteid="1593">
              <RESULTS>
                <RESULT eventid="1111" points="389" reactiontime="+60" swimtime="00:01:27.81" resultid="1594" heatid="3004" lane="2" entrytime="00:01:27.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="411" reactiontime="+91" swimtime="00:00:39.54" resultid="1595" heatid="3048" lane="3" entrytime="00:00:38.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Januszczak" birthdate="2007-02-18" gender="M" nation="POL" license="100515700266" swrid="5198882" athleteid="1527">
              <RESULTS>
                <RESULT eventid="1075" points="386" reactiontime="+68" swimtime="00:00:28.70" resultid="1528" heatid="2968" lane="7" entrytime="00:00:28.48" entrycourse="LCM" />
                <RESULT eventid="1107" points="332" reactiontime="+62" swimtime="00:02:27.20" resultid="1529" heatid="3000" lane="7" entrytime="00:02:25.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:11.05" />
                    <SPLIT distance="150" swimtime="00:01:50.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="276" reactiontime="+54" swimtime="00:00:34.18" resultid="1530" heatid="3021" lane="5" entrytime="00:00:32.15" entrycourse="LCM" />
                <RESULT eventid="1139" points="322" reactiontime="+67" swimtime="00:01:08.38" resultid="1531" heatid="3039" lane="6" entrytime="00:01:03.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Pawlak" birthdate="2005-04-15" gender="M" nation="POL" license="100515700211" swrid="5117073" athleteid="1555">
              <RESULTS>
                <RESULT eventid="1083" points="477" swimtime="00:02:41.32" resultid="1556" heatid="2976" lane="2" entrytime="00:02:38.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                    <SPLIT distance="100" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:57.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="530" reactiontime="+73" swimtime="00:01:10.26" resultid="1557" heatid="3010" lane="9" entrytime="00:01:10.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="545" reactiontime="+70" swimtime="00:00:31.76" resultid="1558" heatid="3057" lane="9" entrytime="00:00:32.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Mazurkiewicz" birthdate="2008-10-03" gender="F" nation="POL" license="100515600299" swrid="5255342" athleteid="1562">
              <RESULTS>
                <RESULT eventid="1087" points="150" reactiontime="+87" swimtime="00:01:44.28" resultid="1563" heatid="2977" lane="4" entrytime="00:01:42.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="159" reactiontime="+77" swimtime="00:00:45.03" resultid="1564" heatid="3013" lane="4" entrytime="00:00:45.31" entrycourse="LCM" />
                <RESULT eventid="1135" points="212" swimtime="00:01:26.69" resultid="1565" heatid="3030" lane="7" entrytime="00:01:22.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Pietrzak" birthdate="2005-03-16" gender="M" nation="POL" license="100515700208" swrid="5117074" athleteid="1509">
              <RESULTS>
                <RESULT eventid="1075" points="468" reactiontime="+75" swimtime="00:00:26.92" resultid="1510" heatid="2969" lane="3" entrytime="00:00:26.76" entrycourse="LCM" />
                <RESULT eventid="1107" points="370" reactiontime="+69" swimtime="00:02:22.03" resultid="1511" heatid="2999" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:08.02" />
                    <SPLIT distance="150" swimtime="00:01:46.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="447" reactiontime="+71" swimtime="00:01:01.35" resultid="1512" heatid="3041" lane="6" entrytime="00:00:58.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Jędrych" birthdate="2004-07-23" gender="M" nation="POL" license="100515700183" swrid="5034201" athleteid="1443">
              <RESULTS>
                <RESULT eventid="1067" points="517" swimtime="00:05:03.81" resultid="1444" heatid="2950" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:08.95" />
                    <SPLIT distance="150" swimtime="00:01:49.04" />
                    <SPLIT distance="200" swimtime="00:02:29.03" />
                    <SPLIT distance="250" swimtime="00:03:11.93" />
                    <SPLIT distance="300" swimtime="00:03:55.89" />
                    <SPLIT distance="350" swimtime="00:04:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="587" reactiontime="+66" swimtime="00:02:01.78" resultid="1445" heatid="3001" lane="4" entrytime="00:02:01.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                    <SPLIT distance="100" swimtime="00:01:00.72" />
                    <SPLIT distance="150" swimtime="00:01:32.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="602" reactiontime="+73" swimtime="00:00:55.55" resultid="1446" heatid="3043" lane="8" entrytime="00:00:55.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="436" reactiontime="+67" swimtime="00:02:30.32" resultid="1447" heatid="3072" lane="7" entrytime="00:02:20.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="150" swimtime="00:01:55.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kornelia" lastname="Kubacka" birthdate="2006-12-16" gender="F" nation="POL" license="100515600254" swrid="4027317" athleteid="1448">
              <RESULTS>
                <RESULT eventid="1071" points="313" reactiontime="+80" swimtime="00:00:34.86" resultid="1449" heatid="2955" lane="8" entrytime="00:00:33.49" entrycourse="LCM" />
                <RESULT eventid="1135" points="263" reactiontime="+78" swimtime="00:01:20.65" resultid="1450" heatid="3031" lane="1" entrytime="00:01:15.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Nowicki" birthdate="1998-08-10" gender="M" nation="POL" license="100515700279" swrid="4711042" athleteid="1500">
              <RESULTS>
                <RESULT eventid="1075" points="462" reactiontime="+79" swimtime="00:00:27.04" resultid="1501" heatid="2963" lane="1" />
                <RESULT eventid="1091" points="476" reactiontime="+74" swimtime="00:01:03.36" resultid="1502" heatid="2982" lane="8" entrytime="00:01:02.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="500" reactiontime="+73" swimtime="00:00:28.04" resultid="1503" heatid="3023" lane="1" entrytime="00:00:27.94" entrycourse="LCM" />
                <RESULT eventid="1171" points="428" reactiontime="+76" swimtime="00:02:31.25" resultid="1504" heatid="3071" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:01:13.04" />
                    <SPLIT distance="150" swimtime="00:01:58.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Brdęk" birthdate="2005-08-23" gender="F" nation="POL" license="100515600221" swrid="5117086" athleteid="1463">
              <RESULTS>
                <RESULT eventid="1071" points="459" reactiontime="+76" swimtime="00:00:30.67" resultid="1464" heatid="2956" lane="3" entrytime="00:00:30.25" entrycourse="LCM" />
                <RESULT eventid="1111" points="475" reactiontime="+76" swimtime="00:01:22.17" resultid="1465" heatid="3004" lane="4" entrytime="00:01:24.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="498" reactiontime="+68" swimtime="00:00:37.08" resultid="1466" heatid="3048" lane="4" entrytime="00:00:37.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Ciszak" birthdate="2006-03-10" gender="F" nation="POL" license="100515600242" swrid="4027104" athleteid="1559">
              <RESULTS>
                <RESULT eventid="1087" points="184" reactiontime="+81" swimtime="00:01:37.48" resultid="1560" heatid="2977" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="240" reactiontime="+86" swimtime="00:03:01.55" resultid="1561" heatid="2994" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:25.97" />
                    <SPLIT distance="150" swimtime="00:02:13.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Brzezicha" birthdate="2008-04-19" gender="M" nation="POL" license="100515700287" swrid="5255303" athleteid="1532">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="1533" heatid="2966" lane="2" entrytime="00:00:31.60" entrycourse="LCM" />
                <RESULT eventid="1115" status="DNS" swimtime="00:00:00.00" resultid="1534" heatid="3008" lane="2" entrytime="00:01:31.94" entrycourse="LCM" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="1535" heatid="3038" lane="3" entrytime="00:01:12.05" entrycourse="LCM" />
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="1536" heatid="3053" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Grzechowiak" birthdate="2006-08-13" gender="M" nation="POL" license="100515700251" swrid="4027106" athleteid="1480">
              <RESULTS>
                <RESULT eventid="1075" points="319" reactiontime="+90" swimtime="00:00:30.59" resultid="1481" heatid="2963" lane="3" />
                <RESULT eventid="1139" points="316" reactiontime="+79" swimtime="00:01:08.87" resultid="1482" heatid="3039" lane="0" entrytime="00:01:07.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Pracharczyk" birthdate="2006-04-05" gender="F" nation="POL" license="100515600243" swrid="4027107" athleteid="1596">
              <RESULTS>
                <RESULT eventid="1127" points="402" reactiontime="+76" swimtime="00:02:47.01" resultid="1597" heatid="3026" lane="6" entrytime="00:02:47.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                    <SPLIT distance="100" swimtime="00:01:20.56" />
                    <SPLIT distance="150" swimtime="00:02:04.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="460" reactiontime="+70" swimtime="00:05:06.26" resultid="1598" heatid="3074" lane="2" entrytime="00:05:07.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:12.34" />
                    <SPLIT distance="150" swimtime="00:01:51.42" />
                    <SPLIT distance="200" swimtime="00:02:30.59" />
                    <SPLIT distance="250" swimtime="00:03:09.98" />
                    <SPLIT distance="300" swimtime="00:03:49.39" />
                    <SPLIT distance="350" swimtime="00:04:29.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymoteusz" lastname="Tomczak" birthdate="2002-05-02" gender="M" nation="POL" license="100515700236" swrid="5071598" athleteid="1551">
              <RESULTS>
                <RESULT eventid="1083" points="613" reactiontime="+67" swimtime="00:02:28.45" resultid="1552" heatid="2976" lane="4" entrytime="00:02:27.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="150" swimtime="00:01:49.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="596" reactiontime="+64" swimtime="00:01:07.56" resultid="1553" heatid="3010" lane="4" entrytime="00:01:06.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="634" reactiontime="+60" swimtime="00:00:30.20" resultid="1554" heatid="3057" lane="5" entrytime="00:00:30.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Bocian" birthdate="2007-07-24" gender="M" nation="POL" license="100515700263" swrid="5198880" athleteid="1522">
              <RESULTS>
                <RESULT eventid="1075" points="349" reactiontime="+76" swimtime="00:00:29.69" resultid="1523" heatid="2967" lane="8" entrytime="00:00:30.07" entrycourse="LCM" />
                <RESULT eventid="1099" points="359" reactiontime="+68" swimtime="00:00:33.74" resultid="1524" heatid="2992" lane="0" entrytime="00:00:33.24" entrycourse="LCM" />
                <RESULT eventid="1123" points="380" reactiontime="+73" swimtime="00:00:30.74" resultid="1525" heatid="3022" lane="0" entrytime="00:00:31.49" entrycourse="LCM" />
                <RESULT eventid="1163" points="350" reactiontime="+77" swimtime="00:01:13.53" resultid="1526" heatid="3064" lane="5" entrytime="00:01:13.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Borys" lastname="Góralczyk" birthdate="2006-04-26" gender="M" nation="POL" license="100515700245" swrid="4951938" athleteid="1483">
              <RESULTS>
                <RESULT eventid="1075" points="376" reactiontime="+99" swimtime="00:00:28.95" resultid="1484" heatid="2960" lane="1" />
                <RESULT eventid="1123" points="344" reactiontime="+70" swimtime="00:00:31.78" resultid="1485" heatid="3019" lane="1" />
                <RESULT eventid="1147" points="334" reactiontime="+70" swimtime="00:00:37.38" resultid="1486" heatid="3054" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Wojtyniak" birthdate="2005-06-16" gender="M" nation="POL" license="100515700217" swrid="5117075" athleteid="1513">
              <RESULTS>
                <RESULT eventid="1075" points="459" reactiontime="+77" swimtime="00:00:27.10" resultid="1514" heatid="2970" lane="9" entrytime="00:00:26.46" entrycourse="LCM" />
                <RESULT eventid="1099" points="435" reactiontime="+58" swimtime="00:00:31.66" resultid="1515" heatid="2992" lane="2" entrytime="00:00:30.30" entrycourse="LCM" />
                <RESULT eventid="1147" points="380" reactiontime="+71" swimtime="00:00:35.82" resultid="1516" heatid="3055" lane="3" entrytime="00:00:39.80" entrycourse="LCM" />
                <RESULT eventid="1163" points="453" reactiontime="+59" swimtime="00:01:07.48" resultid="1517" heatid="3065" lane="7" entrytime="00:01:05.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Depa" birthdate="2004-01-20" gender="M" nation="POL" license="100515700197" swrid="5034193" athleteid="1570">
              <RESULTS>
                <RESULT eventid="1091" points="290" reactiontime="+82" swimtime="00:01:14.78" resultid="1571" heatid="2980" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="481" reactiontime="+72" swimtime="00:02:10.13" resultid="1572" heatid="3000" lane="4" entrytime="00:02:11.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                    <SPLIT distance="100" swimtime="00:01:03.26" />
                    <SPLIT distance="150" swimtime="00:01:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="413" reactiontime="+77" swimtime="00:00:29.89" resultid="1573" heatid="3023" lane="9" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="1139" points="527" reactiontime="+73" swimtime="00:00:58.05" resultid="1574" heatid="3042" lane="9" entrytime="00:00:57.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Apolonia" lastname="Popławska" birthdate="2002-06-01" gender="F" nation="POL" license="100515600277" swrid="4946114" athleteid="1456">
              <RESULTS>
                <RESULT eventid="1071" points="533" reactiontime="+69" swimtime="00:00:29.19" resultid="1457" heatid="2958" lane="6" entrytime="00:00:28.69" entrycourse="LCM" />
                <RESULT eventid="1111" points="462" reactiontime="+73" swimtime="00:01:22.95" resultid="1458" heatid="3005" lane="7" entrytime="00:01:19.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="555" reactiontime="+67" swimtime="00:00:35.76" resultid="1459" heatid="3049" lane="1" entrytime="00:00:35.87" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+64" swimtime="00:01:48.14" resultid="1599" heatid="2948" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.21" />
                    <SPLIT distance="100" swimtime="00:00:50.32" />
                    <SPLIT distance="150" swimtime="00:01:20.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1551" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="1505" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="1460" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="1456" number="4" reactiontime="+2" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1183" reactiontime="+69" swimtime="00:02:01.92" resultid="1601" heatid="3079" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:05.20" />
                    <SPLIT distance="150" swimtime="00:01:31.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1575" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="1456" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="1551" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="1460" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+88" swimtime="00:01:55.16" resultid="1600" heatid="2947" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="100" swimtime="00:00:57.99" />
                    <SPLIT distance="150" swimtime="00:01:28.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1593" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="1589" number="2" />
                    <RELAYPOSITION athleteid="1596" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="1547" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="01" clubid="1602" name="KS Rekin Świebodzice">
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Gajdowska" birthdate="1995-07-17" gender="F" nation="POL" license="102001600173" swrid="4258728" athleteid="1629">
              <RESULTS>
                <RESULT eventid="1071" points="554" reactiontime="+70" swimtime="00:00:28.81" resultid="1630" heatid="2958" lane="4" entrytime="00:00:28.47" entrycourse="LCM" />
                <RESULT eventid="1135" points="591" reactiontime="+66" swimtime="00:01:01.61" resultid="1631" heatid="3034" lane="1" entrytime="00:01:01.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Wajsberg" birthdate="2009-09-29" gender="F" nation="POL" license="102001600154" swrid="5260101" athleteid="1603">
              <RESULTS>
                <RESULT eventid="1071" points="433" reactiontime="+66" swimtime="00:00:31.27" resultid="1604" heatid="2956" lane="1" entrytime="00:00:31.14" entrycourse="LCM" />
                <RESULT eventid="1103" points="388" reactiontime="+77" swimtime="00:02:34.86" resultid="1605" heatid="2995" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:14.04" />
                    <SPLIT distance="150" swimtime="00:01:55.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="401" reactiontime="+69" swimtime="00:01:10.07" resultid="1606" heatid="3031" lane="3" entrytime="00:01:10.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="364" reactiontime="+63" swimtime="00:01:20.59" resultid="1607" heatid="3060" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Brzozowski" birthdate="2006-04-21" gender="M" nation="POL" license="102001700178" swrid="5449489" athleteid="1632">
              <RESULTS>
                <RESULT eventid="1075" points="248" reactiontime="+96" swimtime="00:00:33.27" resultid="1633" heatid="2963" lane="6" />
                <RESULT eventid="1099" points="193" reactiontime="+84" swimtime="00:00:41.51" resultid="1634" heatid="2989" lane="4" />
                <RESULT eventid="1139" points="247" reactiontime="+96" swimtime="00:01:14.75" resultid="1635" heatid="3037" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Folkman" birthdate="2009-10-06" gender="F" nation="POL" license="102001600180" swrid="5449620" athleteid="1624">
              <RESULTS>
                <RESULT eventid="1071" points="323" reactiontime="+91" swimtime="00:00:34.49" resultid="1625" heatid="2955" lane="9" entrytime="00:00:33.87" entrycourse="LCM" />
                <RESULT eventid="1119" points="231" reactiontime="+87" swimtime="00:00:39.78" resultid="1626" heatid="3013" lane="3" />
                <RESULT eventid="1135" points="296" reactiontime="+93" swimtime="00:01:17.53" resultid="1627" heatid="3030" lane="3" entrytime="00:01:20.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="1628" heatid="3067" lane="5" entrytime="00:03:20.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Romanowska" birthdate="2008-10-05" gender="F" nation="POL" license="102001600144" swrid="5263268" athleteid="1612">
              <RESULTS>
                <RESULT eventid="1071" points="364" reactiontime="+93" swimtime="00:00:33.13" resultid="1613" heatid="2952" lane="9" />
                <RESULT eventid="1135" points="349" reactiontime="+89" swimtime="00:01:13.44" resultid="1614" heatid="3031" lane="8" entrytime="00:01:16.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="300" reactiontime="+72" swimtime="00:01:25.98" resultid="1615" heatid="3061" lane="2" entrytime="00:01:27.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Kopeć" birthdate="2008-09-15" gender="M" nation="POL" license="102001700181" swrid="5285302" athleteid="1646">
              <RESULTS>
                <RESULT eventid="1075" points="279" reactiontime="+79" swimtime="00:00:31.98" resultid="1647" heatid="2964" lane="3" />
                <RESULT eventid="1123" points="243" reactiontime="+73" swimtime="00:00:35.67" resultid="1648" heatid="3017" lane="2" />
                <RESULT eventid="1147" points="220" reactiontime="+81" swimtime="00:00:42.95" resultid="1649" heatid="3054" lane="3" />
                <RESULT eventid="1171" points="233" reactiontime="+57" swimtime="00:03:05.12" resultid="1650" heatid="3071" lane="4" entrytime="00:03:00.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:28.56" />
                    <SPLIT distance="150" swimtime="00:02:21.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonina" lastname="Horbacz" birthdate="2007-07-16" gender="F" nation="POL" license="102001600171" swrid="5323392" athleteid="1616">
              <RESULTS>
                <RESULT eventid="1071" points="374" swimtime="00:00:32.84" resultid="1617" heatid="2955" lane="2" entrytime="00:00:32.64" entrycourse="LCM" />
                <RESULT eventid="1119" points="258" reactiontime="+88" swimtime="00:00:38.35" resultid="1618" heatid="3014" lane="8" entrytime="00:00:38.59" entrycourse="LCM" />
                <RESULT eventid="1135" points="338" reactiontime="+71" swimtime="00:01:14.20" resultid="1619" heatid="3031" lane="7" entrytime="00:01:15.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natasza" lastname="Bylińska" birthdate="2007-02-06" gender="F" nation="POL" license="102001600137" swrid="5088581" athleteid="1620">
              <RESULTS>
                <RESULT eventid="1071" points="310" swimtime="00:00:34.94" resultid="1621" heatid="2952" lane="2" />
                <RESULT eventid="1095" points="269" reactiontime="+75" swimtime="00:00:41.77" resultid="1622" heatid="2984" lane="7" />
                <RESULT eventid="1167" points="293" reactiontime="+87" swimtime="00:03:09.80" resultid="1623" heatid="3067" lane="4" entrytime="00:03:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                    <SPLIT distance="100" swimtime="00:01:28.55" />
                    <SPLIT distance="150" swimtime="00:02:27.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aurelia" lastname="Świdurska" birthdate="2009-09-24" gender="F" nation="POL" license="102001600150" swrid="5316783" athleteid="1608">
              <RESULTS>
                <RESULT eventid="1071" points="340" reactiontime="+80" swimtime="00:00:33.91" resultid="1609" heatid="2955" lane="0" entrytime="00:00:33.84" entrycourse="LCM" />
                <RESULT eventid="1135" points="330" reactiontime="+78" swimtime="00:01:14.79" resultid="1610" heatid="3031" lane="0" entrytime="00:01:16.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="332" reactiontime="+78" swimtime="00:03:01.97" resultid="1611" heatid="3068" lane="0" entrytime="00:03:05.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:30.25" />
                    <SPLIT distance="150" swimtime="00:02:21.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Franciszek" lastname="Horbacz" birthdate="2007-07-16" gender="M" nation="POL" license="102001700170" swrid="5260099" athleteid="1641">
              <RESULTS>
                <RESULT eventid="1075" points="318" reactiontime="+66" swimtime="00:00:30.62" resultid="1642" heatid="2967" lane="0" entrytime="00:00:30.19" entrycourse="LCM" />
                <RESULT eventid="1099" points="313" reactiontime="+70" swimtime="00:00:35.33" resultid="1643" heatid="2991" lane="4" entrytime="00:00:34.56" entrycourse="LCM" />
                <RESULT eventid="1123" points="263" reactiontime="+73" swimtime="00:00:34.74" resultid="1644" heatid="3021" lane="2" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1179" points="325" reactiontime="+74" swimtime="00:05:20.02" resultid="1645" heatid="3077" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="150" swimtime="00:01:55.72" />
                    <SPLIT distance="200" swimtime="00:02:37.74" />
                    <SPLIT distance="250" swimtime="00:03:19.45" />
                    <SPLIT distance="300" swimtime="00:04:01.23" />
                    <SPLIT distance="350" swimtime="00:04:42.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Glejzer" birthdate="2006-02-26" gender="M" nation="POL" license="102001700112" swrid="4995330" athleteid="1636">
              <RESULTS>
                <RESULT eventid="1075" points="484" reactiontime="+74" swimtime="00:00:26.62" resultid="1637" heatid="2962" lane="7" />
                <RESULT eventid="1123" points="454" reactiontime="+67" swimtime="00:00:28.97" resultid="1638" heatid="3022" lane="4" entrytime="00:00:29.11" entrycourse="LCM" />
                <RESULT eventid="1139" points="472" swimtime="00:01:00.21" resultid="1639" heatid="3041" lane="2" entrytime="00:00:58.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="439" reactiontime="+72" swimtime="00:02:29.90" resultid="1640" heatid="3069" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:11.22" />
                    <SPLIT distance="150" swimtime="00:01:55.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1183" reactiontime="+69" swimtime="00:02:15.54" resultid="1655" heatid="3079" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                    <SPLIT distance="150" swimtime="00:01:47.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1603" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="1646" number="2" reactiontime="+9" />
                    <RELAYPOSITION athleteid="1636" number="3" />
                    <RELAYPOSITION athleteid="1629" number="4" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="15" clubid="1961" name="KU AZS UAM Poznań">
          <ATHLETES>
            <ATHLETE firstname="Witold" lastname="Świtalski" birthdate="2009-05-09" gender="M" nation="POL" license="103315700051" swrid="5334825" athleteid="1999">
              <RESULTS>
                <RESULT eventid="1075" points="177" reactiontime="+98" swimtime="00:00:37.24" resultid="2000" heatid="2965" lane="3" entrytime="00:00:37.31" entrycourse="LCM" />
                <RESULT eventid="1123" points="139" swimtime="00:00:42.98" resultid="2001" heatid="3021" lane="8" entrytime="00:00:44.98" entrycourse="LCM" />
                <RESULT eventid="1139" points="161" reactiontime="+74" swimtime="00:01:26.17" resultid="2002" heatid="3038" lane="0" entrytime="00:01:25.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matylda" lastname="Ober" birthdate="2008-10-31" gender="F" nation="POL" license="103315600049" swrid="5214664" athleteid="2010">
              <RESULTS>
                <RESULT eventid="1079" points="286" swimtime="00:03:30.90" resultid="2011" heatid="2972" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.79" />
                    <SPLIT distance="100" swimtime="00:01:40.22" />
                    <SPLIT distance="150" swimtime="00:02:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="299" reactiontime="+73" swimtime="00:01:35.86" resultid="2012" heatid="3003" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="311" reactiontime="+80" swimtime="00:00:43.38" resultid="2013" heatid="3047" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olga" lastname="Dolata" birthdate="2008-02-05" gender="F" nation="POL" license="103315600031" swrid="5204346" athleteid="1966">
              <RESULTS>
                <RESULT eventid="1071" points="577" reactiontime="+61" swimtime="00:00:28.43" resultid="1967" heatid="2959" lane="0" entrytime="00:00:28.35" entrycourse="LCM" />
                <RESULT eventid="1103" points="526" reactiontime="+64" swimtime="00:02:19.90" resultid="1968" heatid="2997" lane="1" entrytime="00:02:18.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="100" swimtime="00:01:05.59" />
                    <SPLIT distance="150" swimtime="00:01:43.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="473" reactiontime="+72" swimtime="00:00:37.71" resultid="1969" heatid="3047" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Witold" lastname="Hadyński" birthdate="2010-05-20" gender="M" nation="POL" license="103315700068" swrid="5278394" athleteid="2014">
              <RESULTS>
                <RESULT eventid="1123" points="145" reactiontime="+47" swimtime="00:00:42.36" resultid="2015" heatid="3019" lane="5" />
                <RESULT eventid="1139" points="188" reactiontime="+64" swimtime="00:01:21.76" resultid="2016" heatid="3038" lane="8" entrytime="00:01:20.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olgierd" lastname="Lasik" birthdate="2005-05-09" gender="M" nation="POL" license="103315700024" swrid="5198896" athleteid="1983">
              <RESULTS>
                <RESULT eventid="1075" points="481" reactiontime="+62" swimtime="00:00:26.68" resultid="1984" heatid="2970" lane="0" entrytime="00:00:26.36" entrycourse="LCM" />
                <RESULT eventid="1107" points="460" reactiontime="+71" swimtime="00:02:12.09" resultid="1985" heatid="3001" lane="9" entrytime="00:02:10.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="100" swimtime="00:01:05.09" />
                    <SPLIT distance="150" swimtime="00:01:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="476" swimtime="00:00:33.22" resultid="1986" heatid="3056" lane="2" entrytime="00:00:33.07" entrycourse="LCM" />
                <RESULT eventid="1171" points="481" reactiontime="+61" swimtime="00:02:25.42" resultid="1987" heatid="3072" lane="0" entrytime="00:02:26.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="100" swimtime="00:01:10.35" />
                    <SPLIT distance="150" swimtime="00:01:52.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Cybulski" birthdate="2011-08-26" gender="M" nation="POL" license="103315700091" swrid="5448926" athleteid="2007">
              <RESULTS>
                <RESULT eventid="1075" points="145" reactiontime="+83" swimtime="00:00:39.75" resultid="2008" heatid="2962" lane="1" />
                <RESULT eventid="1139" points="148" swimtime="00:01:28.51" resultid="2009" heatid="3035" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Onichimiuk" birthdate="2008-07-22" gender="F" nation="POL" license="103315600052" swrid="5214734" athleteid="1974">
              <RESULTS>
                <RESULT eventid="1071" points="417" reactiontime="+67" swimtime="00:00:31.68" resultid="1975" heatid="2955" lane="3" entrytime="00:00:32.01" entrycourse="LCM" />
                <RESULT eventid="1119" points="352" swimtime="00:00:34.57" resultid="1976" heatid="3014" lane="7" entrytime="00:00:34.75" entrycourse="LCM" />
                <RESULT eventid="1167" points="414" swimtime="00:02:49.10" resultid="1977" heatid="3067" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:20.67" />
                    <SPLIT distance="150" swimtime="00:02:10.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Kałek" birthdate="2004-01-30" gender="M" nation="POL" license="103315700028" swrid="5198938" athleteid="1978">
              <RESULTS>
                <RESULT eventid="1075" points="383" reactiontime="+66" swimtime="00:00:28.79" resultid="1979" heatid="2968" lane="0" entrytime="00:00:28.85" entrycourse="LCM" />
                <RESULT eventid="1107" points="395" reactiontime="+70" swimtime="00:02:18.97" resultid="1980" heatid="2999" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:07.40" />
                    <SPLIT distance="150" swimtime="00:01:44.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="406" reactiontime="+67" swimtime="00:01:03.30" resultid="1981" heatid="3040" lane="1" entrytime="00:01:02.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="346" reactiontime="+72" swimtime="00:02:42.30" resultid="1982" heatid="3071" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:19.05" />
                    <SPLIT distance="150" swimtime="00:02:05.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Ignatowicz" birthdate="2008-10-10" gender="M" nation="POL" license="103315700168" swrid="5461141" athleteid="1992">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1075" reactiontime="+45" status="DSQ" swimtime="00:00:00.00" resultid="1993" heatid="2966" lane="0" entrytime="00:00:33.48" entrycourse="LCM" />
                <RESULT eventid="1139" points="227" reactiontime="+74" swimtime="00:01:16.88" resultid="1994" heatid="3038" lane="1" entrytime="00:01:15.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antoni" lastname="Pietrzyk" birthdate="2008-10-22" gender="M" nation="POL" license="103315700060" swrid="5311252" athleteid="1988">
              <RESULTS>
                <RESULT eventid="1075" points="328" reactiontime="+64" swimtime="00:00:30.31" resultid="1989" heatid="2966" lane="6" entrytime="00:00:31.34" entrycourse="LCM" />
                <RESULT eventid="1123" points="361" reactiontime="+52" swimtime="00:00:31.27" resultid="1990" heatid="3021" lane="4" entrytime="00:00:31.86" entrycourse="LCM" />
                <RESULT eventid="1171" points="316" reactiontime="+70" swimtime="00:02:47.27" resultid="1991" heatid="3070" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:17.63" />
                    <SPLIT distance="150" swimtime="00:02:09.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Smykowska" birthdate="2006-02-11" gender="F" nation="POL" license="103315600014" swrid="5096901" athleteid="1962">
              <RESULTS>
                <RESULT eventid="1071" points="440" reactiontime="+65" swimtime="00:00:31.11" resultid="1963" heatid="2952" lane="8" />
                <RESULT eventid="1103" status="DNS" swimtime="00:00:00.00" resultid="1964" heatid="2996" lane="3" entrytime="00:02:25.72" entrycourse="LCM" />
                <RESULT eventid="1175" points="437" reactiontime="+67" swimtime="00:05:11.37" resultid="1965" heatid="3073" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:12.81" />
                    <SPLIT distance="150" swimtime="00:01:53.63" />
                    <SPLIT distance="200" swimtime="00:02:34.12" />
                    <SPLIT distance="250" swimtime="00:03:14.28" />
                    <SPLIT distance="300" swimtime="00:03:55.11" />
                    <SPLIT distance="350" swimtime="00:04:34.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konstanty" lastname="Walkowiak" birthdate="2009-04-20" gender="M" nation="POL" license="103315700046" swrid="5214829" athleteid="1995">
              <RESULTS>
                <RESULT eventid="1075" points="200" reactiontime="+49" swimtime="00:00:35.74" resultid="1996" heatid="2965" lane="4" entrytime="00:00:36.16" entrycourse="LCM" />
                <RESULT eventid="1099" points="224" reactiontime="+87" swimtime="00:00:39.49" resultid="1997" heatid="2991" lane="8" entrytime="00:00:37.92" entrycourse="LCM" />
                <RESULT eventid="1163" points="235" reactiontime="+77" swimtime="00:01:23.95" resultid="1998" heatid="3064" lane="1" entrytime="00:01:22.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Wolska" birthdate="2009-01-29" gender="F" nation="POL" athleteid="3080">
              <RESULTS>
                <RESULT eventid="1071" points="267" reactiontime="+88" swimtime="00:00:36.72" resultid="3081" heatid="2951" lane="9" late="yes" />
                <RESULT eventid="1127" points="291" reactiontime="+93" swimtime="00:03:06.03" resultid="3082" heatid="3025" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.98" />
                    <SPLIT distance="100" swimtime="00:01:32.10" />
                    <SPLIT distance="150" swimtime="00:02:20.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="279" reactiontime="+80" swimtime="00:03:12.80" resultid="3083" heatid="3066" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.99" />
                    <SPLIT distance="100" swimtime="00:01:35.18" />
                    <SPLIT distance="150" swimtime="00:02:32.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Kowalik" birthdate="1991-01-05" gender="M" nation="POL" license="103315700017" swrid="4072386" athleteid="2003">
              <RESULTS>
                <RESULT eventid="1075" points="567" reactiontime="+72" swimtime="00:00:25.26" resultid="2004" heatid="2961" lane="8" />
                <RESULT eventid="1099" points="545" reactiontime="+67" swimtime="00:00:29.38" resultid="2005" heatid="2993" lane="1" entrytime="00:00:29.18" entrycourse="LCM" />
                <RESULT eventid="1123" points="604" reactiontime="+63" swimtime="00:00:26.34" resultid="2006" heatid="3024" lane="1" entrytime="00:00:26.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01202" nation="POL" region="02" clubid="1325" name="KP Delfin Inowrocław">
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Kuls" birthdate="2003-04-12" gender="M" nation="POL" license="101202700073" swrid="4827327" athleteid="1330">
              <RESULTS>
                <RESULT eventid="1075" points="574" reactiontime="+72" swimtime="00:00:25.16" resultid="1331" heatid="2971" lane="6" entrytime="00:00:24.74" entrycourse="LCM" />
                <RESULT eventid="1099" points="436" reactiontime="+74" swimtime="00:00:31.64" resultid="1332" heatid="2988" lane="2" />
                <RESULT eventid="1123" points="609" reactiontime="+64" swimtime="00:00:26.27" resultid="1333" heatid="3024" lane="2" entrytime="00:00:25.90" entrycourse="LCM" />
                <RESULT eventid="1147" points="518" reactiontime="+76" swimtime="00:00:32.31" resultid="1334" heatid="3051" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Suchodolski" birthdate="2004-05-12" gender="M" nation="POL" license="101202700098" swrid="5120317" athleteid="1335">
              <RESULTS>
                <RESULT eventid="1083" points="466" reactiontime="+84" swimtime="00:02:42.64" resultid="1336" heatid="2975" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:16.54" />
                    <SPLIT distance="150" swimtime="00:01:59.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="446" reactiontime="+71" swimtime="00:01:14.44" resultid="1337" heatid="3009" lane="1" entrytime="00:01:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="452" reactiontime="+78" swimtime="00:02:28.54" resultid="1338" heatid="3071" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                    <SPLIT distance="100" swimtime="00:01:09.86" />
                    <SPLIT distance="150" swimtime="00:01:52.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Meyer" birthdate="2002-12-10" gender="M" nation="POL" license="101202700116" swrid="5411140" athleteid="1326">
              <RESULTS>
                <RESULT eventid="1075" points="546" reactiontime="+68" swimtime="00:00:25.57" resultid="1327" heatid="2971" lane="0" entrytime="00:00:25.05" entrycourse="LCM" />
                <RESULT eventid="1123" points="573" reactiontime="+83" swimtime="00:00:26.80" resultid="1328" heatid="3019" lane="8" />
                <RESULT eventid="1139" points="555" reactiontime="+70" swimtime="00:00:57.06" resultid="1329" heatid="3042" lane="2" entrytime="00:00:56.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03015" nation="POL" region="15" clubid="2587" name="UKS Fala Swarzędz">
          <ATHLETES>
            <ATHLETE firstname="Oskar" lastname="Szymański" birthdate="2003-08-16" gender="M" nation="POL" license="103015700027" swrid="4947381" athleteid="2608">
              <RESULTS>
                <RESULT eventid="1075" points="467" swimtime="00:00:26.95" resultid="2609" heatid="2969" lane="2" entrytime="00:00:26.95" entrycourse="LCM" />
                <RESULT eventid="1115" points="334" swimtime="00:01:21.91" resultid="2610" heatid="3007" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="386" reactiontime="+64" swimtime="00:00:30.56" resultid="2611" heatid="3018" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Różańska" birthdate="2011-08-13" gender="F" nation="POL" license="103015600060" swrid="5448039" athleteid="2588">
              <RESULTS>
                <RESULT eventid="1071" points="163" reactiontime="+51" swimtime="00:00:43.33" resultid="2589" heatid="2951" lane="6" />
                <RESULT eventid="1143" points="147" swimtime="00:00:55.65" resultid="2590" heatid="3045" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymon" lastname="Waligóra" birthdate="2008-04-03" gender="M" nation="POL" license="103015700039" swrid="4981604" athleteid="2624">
              <RESULTS>
                <RESULT eventid="1083" points="243" reactiontime="+72" swimtime="00:03:21.85" resultid="2625" heatid="2974" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                    <SPLIT distance="100" swimtime="00:01:34.94" />
                    <SPLIT distance="150" swimtime="00:02:29.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="245" reactiontime="+56" swimtime="00:00:41.45" resultid="2626" heatid="3055" lane="7" entrytime="00:00:41.22" entrycourse="LCM" />
                <RESULT eventid="1171" points="185" reactiontime="+65" swimtime="00:03:19.76" resultid="2627" heatid="3070" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:37.83" />
                    <SPLIT distance="150" swimtime="00:02:33.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lea" lastname="Różańska" birthdate="2009-04-30" gender="F" nation="POL" license="103015600045" swrid="5325107" athleteid="2620">
              <RESULTS>
                <RESULT eventid="1079" points="300" reactiontime="+83" swimtime="00:03:27.62" resultid="2621" heatid="2972" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                    <SPLIT distance="100" swimtime="00:01:39.37" />
                    <SPLIT distance="150" swimtime="00:02:33.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="295" reactiontime="+67" swimtime="00:01:36.31" resultid="2622" heatid="3002" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="283" reactiontime="+78" swimtime="00:03:12.08" resultid="2623" heatid="3066" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:31.51" />
                    <SPLIT distance="150" swimtime="00:02:26.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Szmyt" birthdate="2003-04-16" gender="M" nation="POL" license="103015700022" swrid="4920334" athleteid="2591">
              <RESULTS>
                <RESULT eventid="1075" points="557" reactiontime="+79" swimtime="00:00:25.41" resultid="2592" heatid="2971" lane="9" entrytime="00:00:25.12" entrycourse="LCM" />
                <RESULT eventid="1099" points="606" reactiontime="+72" swimtime="00:00:28.35" resultid="2593" heatid="2993" lane="3" entrytime="00:00:28.43" entrycourse="LCM" />
                <RESULT eventid="1139" points="629" reactiontime="+73" swimtime="00:00:54.74" resultid="2594" heatid="3036" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="564" reactiontime="+78" swimtime="00:01:02.75" resultid="2595" heatid="3063" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Adamczyk" birthdate="2005-03-04" gender="M" nation="POL" license="103015700032" swrid="5179131" athleteid="2604">
              <RESULTS>
                <RESULT eventid="1075" points="476" reactiontime="+73" swimtime="00:00:26.78" resultid="2605" heatid="2969" lane="7" entrytime="00:00:27.17" entrycourse="LCM" />
                <RESULT eventid="1107" points="420" reactiontime="+76" swimtime="00:02:16.12" resultid="2606" heatid="2999" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="100" swimtime="00:01:05.78" />
                    <SPLIT distance="150" swimtime="00:01:41.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="500" reactiontime="+64" swimtime="00:00:59.09" resultid="2607" heatid="3040" lane="4" entrytime="00:01:00.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Waligóra" birthdate="2006-01-28" gender="M" nation="POL" license="103015700038" swrid="5179132" athleteid="2612">
              <RESULTS>
                <RESULT eventid="1075" points="468" reactiontime="+79" swimtime="00:00:26.92" resultid="2613" heatid="2969" lane="9" entrytime="00:00:27.53" entrycourse="LCM" />
                <RESULT eventid="1123" points="475" reactiontime="+71" swimtime="00:00:28.54" resultid="2614" heatid="3022" lane="3" entrytime="00:00:29.36" entrycourse="LCM" />
                <RESULT eventid="1139" points="503" reactiontime="+67" swimtime="00:00:58.95" resultid="2615" heatid="3040" lane="5" entrytime="00:01:00.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="420" reactiontime="+69" swimtime="00:04:53.73" resultid="2616" heatid="3076" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="100" swimtime="00:01:07.40" />
                    <SPLIT distance="150" swimtime="00:01:44.76" />
                    <SPLIT distance="200" swimtime="00:02:22.60" />
                    <SPLIT distance="250" swimtime="00:03:01.74" />
                    <SPLIT distance="300" swimtime="00:03:40.68" />
                    <SPLIT distance="350" swimtime="00:04:19.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksy" lastname="Bielawski" birthdate="2009-04-24" gender="M" nation="POL" license="103015700074" swrid="5461132" athleteid="2617">
              <RESULTS>
                <RESULT eventid="1075" points="254" reactiontime="+56" swimtime="00:00:33.01" resultid="2618" heatid="2966" lane="9" entrytime="00:00:34.68" entrycourse="LCM" />
                <RESULT eventid="1139" points="206" reactiontime="+63" swimtime="00:01:19.38" resultid="2619" heatid="3038" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Wermiński" birthdate="2004-09-26" gender="M" nation="POL" license="103015700016" swrid="5096951" athleteid="2596">
              <RESULTS>
                <RESULT eventid="1075" points="561" reactiontime="+79" swimtime="00:00:25.34" resultid="2597" heatid="2970" lane="3" entrytime="00:00:25.51" entrycourse="LCM" />
                <RESULT eventid="1115" points="601" reactiontime="+71" swimtime="00:01:07.37" resultid="2598" heatid="3010" lane="6" entrytime="00:01:08.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="648" reactiontime="+87" swimtime="00:00:29.98" resultid="2599" heatid="3057" lane="4" entrytime="00:00:30.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Marszałkiewicz" birthdate="2003-10-31" gender="M" nation="POL" license="103015700029" swrid="5202983" athleteid="2600">
              <RESULTS>
                <RESULT eventid="1075" points="441" reactiontime="+66" swimtime="00:00:27.46" resultid="2601" heatid="2969" lane="5" entrytime="00:00:26.74" entrycourse="LCM" />
                <RESULT eventid="1107" points="388" reactiontime="+82" swimtime="00:02:19.76" resultid="2602" heatid="2998" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:43.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="458" reactiontime="+71" swimtime="00:00:28.89" resultid="2603" heatid="3023" lane="0" entrytime="00:00:28.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antoni" lastname="Zawadka" birthdate="2008-05-28" gender="M" nation="POL" license="103015700058" swrid="5405704" athleteid="2628">
              <RESULTS>
                <RESULT eventid="1091" points="145" reactiontime="+67" swimtime="00:01:34.18" resultid="2629" heatid="2980" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="230" reactiontime="+48" swimtime="00:00:36.33" resultid="2630" heatid="3019" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00309" nation="POL" region="09" clubid="2141" name="MKS Juvenia Białystok">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Żmiejko" birthdate="1963-01-16" gender="M" nation="POL" license="500309700377" swrid="4186249" athleteid="2142">
              <RESULTS>
                <RESULT eventid="1075" points="361" reactiontime="+88" swimtime="00:00:29.35" resultid="2143" heatid="2964" lane="7" />
                <RESULT eventid="1123" points="367" reactiontime="+87" swimtime="00:00:31.10" resultid="2144" heatid="3018" lane="8" />
                <RESULT eventid="1139" points="361" reactiontime="+87" swimtime="00:01:05.83" resultid="2145" heatid="3037" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03415" nation="POL" region="15" clubid="2488" name="Uks Cityzen">
          <ATHLETES>
            <ATHLETE firstname="Sławomir" lastname="Cybertowicz" birthdate="1966-01-12" gender="M" nation="POL" license="503415700177" swrid="4269915" athleteid="2581">
              <RESULTS>
                <RESULT eventid="1115" points="283" reactiontime="+77" swimtime="00:01:26.57" resultid="2582" heatid="3007" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="303" reactiontime="+67" swimtime="00:00:38.62" resultid="2583" heatid="3053" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alex" lastname="Baranowski" birthdate="2007-02-27" gender="M" nation="POL" license="103415700115" swrid="5405709" athleteid="2513">
              <RESULTS>
                <RESULT eventid="1075" points="410" reactiontime="+79" swimtime="00:00:28.13" resultid="2514" heatid="2961" lane="9" />
                <RESULT eventid="1123" points="352" reactiontime="+72" swimtime="00:00:31.52" resultid="2515" heatid="3021" lane="3" entrytime="00:00:32.59" entrycourse="LCM" />
                <RESULT eventid="1139" points="454" swimtime="00:01:01.00" resultid="2516" heatid="3040" lane="2" entrytime="00:01:01.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Łoboda" birthdate="2008-04-09" gender="F" nation="POL" license="103415600107" swrid="5154973" athleteid="2563">
              <RESULTS>
                <RESULT eventid="1103" points="453" reactiontime="+74" swimtime="00:02:27.09" resultid="2564" heatid="2995" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                    <SPLIT distance="150" swimtime="00:01:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="394" reactiontime="+64" swimtime="00:00:33.30" resultid="2565" heatid="3012" lane="4" />
                <RESULT eventid="1143" points="379" reactiontime="+71" swimtime="00:00:40.60" resultid="2566" heatid="3046" lane="7" />
                <RESULT eventid="1159" points="421" reactiontime="+67" swimtime="00:01:16.79" resultid="2567" heatid="3061" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Liberski" birthdate="2007-05-02" gender="M" nation="POL" license="103415700045" swrid="5096972" athleteid="2522">
              <RESULTS>
                <RESULT eventid="1075" points="381" reactiontime="+67" swimtime="00:00:28.83" resultid="2523" heatid="2960" lane="7" />
                <RESULT eventid="1123" points="352" reactiontime="+64" swimtime="00:00:31.52" resultid="2524" heatid="3019" lane="2" />
                <RESULT eventid="1139" points="418" reactiontime="+69" swimtime="00:01:02.70" resultid="2525" heatid="3037" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Boryski" birthdate="1951-03-05" gender="M" nation="POL" license="503415700180" swrid="4754708" athleteid="2553">
              <RESULTS>
                <RESULT eventid="1099" points="146" reactiontime="+100" swimtime="00:00:45.56" resultid="2554" heatid="2989" lane="9" />
                <RESULT eventid="1131" points="110" reactiontime="+92" swimtime="00:03:53.23" resultid="2555" heatid="3028" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.23" />
                    <SPLIT distance="100" swimtime="00:01:56.45" />
                    <SPLIT distance="150" swimtime="00:02:57.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="109" reactiontime="+112" swimtime="00:07:39.91" resultid="2556" heatid="3077" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.30" />
                    <SPLIT distance="100" swimtime="00:01:51.65" />
                    <SPLIT distance="150" swimtime="00:02:51.03" />
                    <SPLIT distance="200" swimtime="00:03:48.78" />
                    <SPLIT distance="250" swimtime="00:04:47.85" />
                    <SPLIT distance="300" swimtime="00:05:45.56" />
                    <SPLIT distance="350" swimtime="00:06:44.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kostiantyn" lastname="Surkov" birthdate="2006-07-05" gender="M" nation="POL" license="103415700088" swrid="5058525" athleteid="2517">
              <RESULTS>
                <RESULT eventid="1075" points="299" reactiontime="+73" swimtime="00:00:31.24" resultid="2518" heatid="2966" lane="7" entrytime="00:00:31.77" entrycourse="LCM" />
                <RESULT eventid="1115" points="266" reactiontime="+66" swimtime="00:01:28.39" resultid="2519" heatid="3008" lane="6" entrytime="00:01:27.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="340" reactiontime="+73" swimtime="00:01:07.18" resultid="2520" heatid="3038" lane="4" entrytime="00:01:10.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="261" reactiontime="+62" swimtime="00:00:40.56" resultid="2521" heatid="3054" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Gulczyńska" birthdate="2007-08-25" gender="F" nation="POL" license="103415600093" swrid="5198895" athleteid="2489">
              <RESULTS>
                <RESULT eventid="1071" points="547" reactiontime="+69" swimtime="00:00:28.93" resultid="2490" heatid="2956" lane="6" entrytime="00:00:30.33" entrycourse="LCM" />
                <RESULT eventid="1119" points="435" reactiontime="+74" swimtime="00:00:32.23" resultid="2491" heatid="3015" lane="9" entrytime="00:00:32.95" entrycourse="LCM" />
                <RESULT eventid="1143" points="496" reactiontime="+70" swimtime="00:00:37.14" resultid="2492" heatid="3049" lane="9" entrytime="00:00:37.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Gorzeń" birthdate="2003-01-20" gender="F" nation="POL" license="103415600013" swrid="5071599" athleteid="2500">
              <RESULTS>
                <RESULT eventid="1071" points="454" reactiontime="+73" swimtime="00:00:30.78" resultid="2501" heatid="2953" lane="8" />
                <RESULT eventid="1095" points="454" reactiontime="+76" swimtime="00:00:35.08" resultid="2502" heatid="2983" lane="3" />
                <RESULT eventid="1135" points="446" reactiontime="+53" swimtime="00:01:07.64" resultid="2503" heatid="3029" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kaczmarek" birthdate="1982-10-03" gender="M" nation="POL" license="503415700331" athleteid="2504">
              <RESULTS>
                <RESULT eventid="1075" points="356" reactiontime="+91" swimtime="00:00:29.48" resultid="2505" heatid="2964" lane="6" />
                <RESULT eventid="1083" points="293" reactiontime="+112" swimtime="00:03:09.87" resultid="2506" heatid="2974" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.48" />
                    <SPLIT distance="100" swimtime="00:01:30.16" />
                    <SPLIT distance="150" swimtime="00:02:20.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="284" reactiontime="+96" swimtime="00:01:26.46" resultid="2507" heatid="3007" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="340" reactiontime="+100" swimtime="00:01:07.21" resultid="2508" heatid="3037" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Łutowicz" birthdate="1950-08-23" gender="F" nation="POL" license="503415600183" swrid="4188428" athleteid="2493">
              <RESULTS>
                <RESULT eventid="1071" points="162" reactiontime="+98" swimtime="00:00:43.39" resultid="2494" heatid="2952" lane="3" />
                <RESULT eventid="1119" points="76" reactiontime="+100" swimtime="00:00:57.67" resultid="2495" heatid="3013" lane="0" />
                <RESULT eventid="1159" points="99" reactiontime="+92" swimtime="00:02:04.31" resultid="2496" heatid="3061" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Pupka" birthdate="2004-05-02" gender="M" nation="POL" license="103415700057" swrid="4981596" athleteid="2571">
              <RESULTS>
                <RESULT eventid="1107" points="429" reactiontime="+78" swimtime="00:02:15.21" resultid="2572" heatid="2998" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:06.26" />
                    <SPLIT distance="150" swimtime="00:01:41.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="486" reactiontime="+66" swimtime="00:04:39.73" resultid="2573" heatid="3076" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:06.83" />
                    <SPLIT distance="150" swimtime="00:01:42.47" />
                    <SPLIT distance="200" swimtime="00:02:18.37" />
                    <SPLIT distance="250" swimtime="00:02:54.05" />
                    <SPLIT distance="300" swimtime="00:03:29.77" />
                    <SPLIT distance="350" swimtime="00:04:05.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Koprowski" birthdate="2003-07-11" gender="M" nation="POL" license="103415700065" swrid="4981652" athleteid="2509">
              <RESULTS>
                <RESULT eventid="1075" points="473" reactiontime="+80" swimtime="00:00:26.82" resultid="2510" heatid="2962" lane="3" />
                <RESULT eventid="1107" points="542" reactiontime="+81" swimtime="00:02:05.10" resultid="2511" heatid="2999" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="100" swimtime="00:01:00.03" />
                    <SPLIT distance="150" swimtime="00:01:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="535" reactiontime="+70" swimtime="00:00:57.75" resultid="2512" heatid="3036" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Bosiacki" birthdate="2007-01-22" gender="M" nation="POL" license="103415700068" swrid="5278372" athleteid="2545">
              <RESULTS>
                <RESULT eventid="1099" points="295" reactiontime="+72" swimtime="00:00:36.04" resultid="2546" heatid="2989" lane="3" />
                <RESULT eventid="1139" points="321" reactiontime="+75" swimtime="00:01:08.49" resultid="2547" heatid="3039" lane="9" entrytime="00:01:10.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="346" reactiontime="+73" swimtime="00:00:36.94" resultid="2548" heatid="3056" lane="0" entrytime="00:00:36.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Pietraszewski" birthdate="1955-04-07" gender="M" nation="POL" license="503415700182" swrid="4187282" athleteid="2584">
              <RESULTS>
                <RESULT eventid="1131" points="163" reactiontime="+89" swimtime="00:03:24.70" resultid="2585" heatid="3028" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.20" />
                    <SPLIT distance="100" swimtime="00:01:39.92" />
                    <SPLIT distance="150" swimtime="00:02:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="159" reactiontime="+93" swimtime="00:01:35.51" resultid="2586" heatid="3063" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Norbert" lastname="Gorzeń" birthdate="2006-06-03" gender="M" nation="POL" license="103415700019" swrid="5138790" athleteid="2534">
              <RESULTS>
                <RESULT eventid="1075" points="387" reactiontime="+81" swimtime="00:00:28.68" resultid="2535" heatid="2964" lane="5" />
                <RESULT eventid="1107" points="412" reactiontime="+72" swimtime="00:02:16.99" resultid="2536" heatid="3000" lane="3" entrytime="00:02:17.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:05.80" />
                    <SPLIT distance="150" swimtime="00:01:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="433" reactiontime="+77" swimtime="00:04:50.89" resultid="2537" heatid="3077" lane="1" entrytime="00:04:58.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                    <SPLIT distance="100" swimtime="00:01:09.74" />
                    <SPLIT distance="150" swimtime="00:01:47.08" />
                    <SPLIT distance="200" swimtime="00:02:24.11" />
                    <SPLIT distance="250" swimtime="00:03:00.73" />
                    <SPLIT distance="300" swimtime="00:03:37.70" />
                    <SPLIT distance="350" swimtime="00:04:15.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Głuszkowski" birthdate="2001-09-24" gender="M" nation="POL" license="103415700008" swrid="4586995" athleteid="2568">
              <RESULTS>
                <RESULT eventid="1179" points="650" reactiontime="+64" swimtime="00:04:13.96" resultid="2570" heatid="3077" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                    <SPLIT distance="100" swimtime="00:01:00.06" />
                    <SPLIT distance="150" swimtime="00:01:31.81" />
                    <SPLIT distance="200" swimtime="00:02:04.28" />
                    <SPLIT distance="250" swimtime="00:02:36.54" />
                    <SPLIT distance="300" swimtime="00:03:09.23" />
                    <SPLIT distance="350" swimtime="00:03:41.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Nochowicz" birthdate="1951-06-03" gender="M" nation="POL" license="503415700186" athleteid="2557">
              <RESULTS>
                <RESULT eventid="1099" points="71" reactiontime="+98" swimtime="00:00:57.94" resultid="2558" heatid="2988" lane="7" />
                <RESULT eventid="1123" points="56" reactiontime="+123" swimtime="00:00:58.05" resultid="2559" heatid="3019" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teresa" lastname="Barełkowska" birthdate="1948-08-02" gender="F" nation="POL" license="503415600350" swrid="4920301" athleteid="2542">
              <RESULTS>
                <RESULT eventid="1095" points="49" reactiontime="+89" swimtime="00:01:13.46" resultid="2543" heatid="2984" lane="1" />
                <RESULT eventid="1143" points="70" swimtime="00:01:11.28" resultid="2544" heatid="3046" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Troszczyński" birthdate="2007-12-16" gender="M" nation="POL" license="103415700094" swrid="5198889" athleteid="2538">
              <RESULTS>
                <RESULT eventid="1091" points="416" reactiontime="+71" swimtime="00:01:06.29" resultid="2539" heatid="2981" lane="3" entrytime="00:01:08.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="383" reactiontime="+76" swimtime="00:00:33.02" resultid="2540" heatid="2992" lane="8" entrytime="00:00:32.36" entrycourse="LCM" />
                <RESULT eventid="1123" points="381" reactiontime="+74" swimtime="00:00:30.71" resultid="2541" heatid="3022" lane="7" entrytime="00:00:30.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Majak" birthdate="2005-07-27" gender="M" nation="POL" license="103415700022" swrid="5096949" athleteid="2574">
              <RESULTS>
                <RESULT eventid="1107" points="351" reactiontime="+80" swimtime="00:02:24.47" resultid="2575" heatid="2998" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:09.38" />
                    <SPLIT distance="150" swimtime="00:01:47.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="395" reactiontime="+75" swimtime="00:04:59.91" resultid="2576" heatid="3075" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:09.45" />
                    <SPLIT distance="150" swimtime="00:01:48.54" />
                    <SPLIT distance="200" swimtime="00:02:27.16" />
                    <SPLIT distance="250" swimtime="00:03:06.41" />
                    <SPLIT distance="300" swimtime="00:03:44.81" />
                    <SPLIT distance="350" swimtime="00:04:23.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Barczyk" birthdate="2007-01-07" gender="M" nation="POL" license="103415700062" swrid="5004223" athleteid="2530">
              <RESULTS>
                <RESULT eventid="1075" points="398" reactiontime="+86" swimtime="00:00:28.42" resultid="2531" heatid="2965" lane="8" />
                <RESULT eventid="1099" points="372" reactiontime="+72" swimtime="00:00:33.37" resultid="2532" heatid="2990" lane="1" />
                <RESULT eventid="1123" points="362" reactiontime="+71" swimtime="00:00:31.23" resultid="2533" heatid="3017" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Miśkiewicz" birthdate="1959-03-24" gender="M" nation="POL" license="503415700185" swrid="4920302" athleteid="2560">
              <RESULTS>
                <RESULT eventid="1099" points="128" reactiontime="+88" swimtime="00:00:47.55" resultid="2561" heatid="2989" lane="8" />
                <RESULT eventid="1163" points="113" reactiontime="+95" swimtime="00:01:47.01" resultid="2562" heatid="3063" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Kaczmarek" birthdate="2007-12-22" gender="M" nation="POL" license="103415700092" swrid="5198919" athleteid="2549">
              <RESULTS>
                <RESULT eventid="1099" points="464" reactiontime="+63" swimtime="00:00:30.99" resultid="2550" heatid="2992" lane="7" entrytime="00:00:31.54" entrycourse="LCM" />
                <RESULT eventid="1147" points="393" reactiontime="+63" swimtime="00:00:35.41" resultid="2551" heatid="3054" lane="1" />
                <RESULT eventid="1163" points="489" reactiontime="+57" swimtime="00:01:05.80" resultid="2552" heatid="3065" lane="8" entrytime="00:01:06.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Łasińska-Błachowicz" birthdate="1954-07-13" gender="F" nation="POL" license="503415600184" athleteid="2497">
              <RESULTS>
                <RESULT eventid="1071" points="101" reactiontime="+111" swimtime="00:00:50.75" resultid="2498" heatid="2953" lane="4" />
                <RESULT eventid="1119" points="64" reactiontime="+127" swimtime="00:01:00.82" resultid="2499" heatid="3013" lane="8" />
                <RESULT eventid="1159" points="70" reactiontime="+102" swimtime="00:02:19.52" resultid="2946" heatid="3061" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Jarzina" birthdate="2007-11-11" gender="M" nation="POL" license="103415700056" swrid="5297966" athleteid="2526">
              <RESULTS>
                <RESULT eventid="1075" points="264" reactiontime="+77" swimtime="00:00:32.58" resultid="2527" heatid="2961" lane="7" />
                <RESULT eventid="1139" points="271" reactiontime="+76" swimtime="00:01:12.43" resultid="2528" heatid="3037" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="199" reactiontime="+76" swimtime="00:00:44.39" resultid="2529" heatid="3050" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Matyszczak" birthdate="1970-12-14" gender="M" nation="POL" license="503415700353" athleteid="2577">
              <RESULTS>
                <RESULT eventid="1107" points="209" reactiontime="+96" swimtime="00:02:51.85" resultid="2578" heatid="2998" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="150" swimtime="00:02:03.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="271" reactiontime="+82" swimtime="00:01:12.45" resultid="2579" heatid="3035" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="168" reactiontime="+96" swimtime="00:01:33.86" resultid="2580" heatid="3063" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="307" reactiontime="+95" swimtime="00:00:30.99" resultid="2945" heatid="2960" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06301" nation="POL" region="01" clubid="2636" name="UKS RAPID Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Oskar" lastname="Gołębiowski" birthdate="2011-03-22" gender="M" nation="POL" license="106301700065" swrid="5450893" athleteid="2642">
              <RESULTS>
                <RESULT eventid="1075" points="62" swimtime="00:00:52.70" resultid="2643" heatid="2965" lane="1" entrytime="00:00:50.58" entrycourse="LCM" />
                <RESULT eventid="1147" points="69" swimtime="00:01:03.24" resultid="2644" heatid="3055" lane="9" entrytime="00:01:05.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Gołębiowski" birthdate="2009-03-03" gender="M" nation="POL" license="106301700030" swrid="5418459" athleteid="2645">
              <RESULTS>
                <RESULT eventid="1083" points="206" swimtime="00:03:33.26" resultid="2646" heatid="2975" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.17" />
                    <SPLIT distance="100" swimtime="00:01:43.88" />
                    <SPLIT distance="150" swimtime="00:02:39.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="171" reactiontime="+60" swimtime="00:01:42.31" resultid="2647" heatid="3007" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="144" reactiontime="+66" swimtime="00:00:49.44" resultid="2648" heatid="3055" lane="0" entrytime="00:00:49.92" entrycourse="LCM" />
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /M10" eventid="1171" reactiontime="+63" status="DSQ" swimtime="00:00:00.00" resultid="2649" heatid="3071" lane="3" entrytime="00:03:19.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.86" />
                    <SPLIT distance="100" swimtime="00:01:45.08" />
                    <SPLIT distance="150" swimtime="00:02:39.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Barczewska" birthdate="2008-09-05" gender="F" nation="POL" license="106301600021" swrid="5418461" athleteid="2637">
              <RESULTS>
                <RESULT eventid="1071" points="261" reactiontime="+85" swimtime="00:00:37.00" resultid="2638" heatid="2954" lane="1" entrytime="00:00:37.67" entrycourse="LCM" />
                <RESULT eventid="1111" points="217" reactiontime="+84" swimtime="00:01:46.67" resultid="2639" heatid="3003" lane="4" entrytime="00:01:44.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="197" reactiontime="+70" swimtime="00:01:28.74" resultid="2640" heatid="3030" lane="1" entrytime="00:01:23.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="210" reactiontime="+83" swimtime="00:00:49.46" resultid="2641" heatid="3046" lane="0" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01610" nation="POL" region="10" clubid="1262" name="Grupa Pływacka Gdynia Masters">
          <ATHLETES>
            <ATHLETE firstname="Czesław" lastname="Mikołajczyk" birthdate="1950-05-18" gender="M" nation="POL" license="501610700006" swrid="4754640" athleteid="1267">
              <RESULTS>
                <RESULT eventid="1083" points="81" reactiontime="+115" swimtime="00:04:50.62" resultid="1268" heatid="2975" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.88" />
                    <SPLIT distance="100" swimtime="00:02:21.02" />
                    <SPLIT distance="150" swimtime="00:03:36.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="76" reactiontime="+112" swimtime="00:02:14.16" resultid="1269" heatid="3006" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="99" reactiontime="+111" swimtime="00:00:56.03" resultid="1270" heatid="3054" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Jacaszek" birthdate="1953-01-24" gender="M" nation="POL" license="501610700018" swrid="4992743" athleteid="1263">
              <RESULTS>
                <RESULT eventid="1083" points="148" reactiontime="+113" swimtime="00:03:58.09" resultid="1264" heatid="2975" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.67" />
                    <SPLIT distance="100" swimtime="00:01:54.44" />
                    <SPLIT distance="150" swimtime="00:02:58.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="167" reactiontime="+107" swimtime="00:01:43.10" resultid="1265" heatid="3006" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="207" reactiontime="+96" swimtime="00:00:43.85" resultid="1266" heatid="3054" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ryszard" lastname="Wachowski" birthdate="1969-09-07" gender="M" nation="POL" license="501610700047" athleteid="1271">
              <RESULTS>
                <RESULT eventid="1123" points="274" reactiontime="+88" swimtime="00:00:34.26" resultid="1272" heatid="3020" lane="2" />
                <RESULT eventid="1171" points="227" reactiontime="+87" swimtime="00:03:06.72" resultid="1273" heatid="3071" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                    <SPLIT distance="150" swimtime="00:02:21.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00704" nation="POL" region="04" clubid="1280" name="Klub Pływacki STILON Gorzów Wlkp.">
          <ATHLETES>
            <ATHLETE firstname="Maksymilian" lastname="Wałcerz" birthdate="2004-07-07" gender="M" nation="POL" license="100704700020" swrid="5084094" athleteid="1293">
              <RESULTS>
                <RESULT eventid="1075" points="581" reactiontime="+77" swimtime="00:00:25.05" resultid="1294" heatid="2971" lane="2" entrytime="00:00:24.80" entrycourse="LCM" />
                <RESULT eventid="1099" points="553" reactiontime="+69" swimtime="00:00:29.23" resultid="1295" heatid="2993" lane="6" entrytime="00:00:28.95" entrycourse="LCM" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="1296" heatid="3043" lane="7" entrytime="00:00:55.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Seń" birthdate="2005-01-28" gender="M" nation="POL" license="100704700018" swrid="5084088" athleteid="1297">
              <RESULTS>
                <RESULT eventid="1091" points="451" reactiontime="+70" swimtime="00:01:04.54" resultid="1298" heatid="2981" lane="4" entrytime="00:01:05.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="371" reactiontime="+66" swimtime="00:01:19.11" resultid="1299" heatid="3008" lane="4" entrytime="00:01:18.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="1300" heatid="3056" lane="8" entrytime="00:00:34.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nikola" lastname="Chorąziak" birthdate="2006-02-21" gender="F" nation="POL" license="100704600041" swrid="5101129" athleteid="1281">
              <RESULTS>
                <RESULT eventid="1071" points="388" reactiontime="+68" swimtime="00:00:32.44" resultid="1282" heatid="2955" lane="6" entrytime="00:00:32.32" entrycourse="LCM" />
                <RESULT eventid="1119" points="344" reactiontime="+66" swimtime="00:00:34.86" resultid="1283" heatid="3014" lane="6" entrytime="00:00:34.40" entrycourse="LCM" />
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="1284" heatid="3048" lane="8" entrytime="00:00:40.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Lech" birthdate="2006-09-24" gender="M" nation="POL" license="100704700032" swrid="4132745" athleteid="1285">
              <RESULTS>
                <RESULT eventid="1075" points="438" reactiontime="+82" swimtime="00:00:27.52" resultid="1286" heatid="2969" lane="1" entrytime="00:00:27.22" entrycourse="LCM" />
                <RESULT eventid="1123" points="341" reactiontime="+83" swimtime="00:00:31.85" resultid="1287" heatid="3022" lane="8" entrytime="00:00:31.49" entrycourse="LCM" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="1288" heatid="3040" lane="3" entrytime="00:01:00.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Kaczmarczyk" birthdate="2003-05-30" gender="M" nation="POL" license="100704700022" swrid="5011820" athleteid="1289">
              <RESULTS>
                <RESULT eventid="1075" points="471" reactiontime="+87" swimtime="00:00:26.86" resultid="1290" heatid="2965" lane="5" entrytime="00:00:37.05" entrycourse="LCM" />
                <RESULT eventid="1091" points="483" reactiontime="+74" swimtime="00:01:03.06" resultid="1291" heatid="2982" lane="0" entrytime="00:01:02.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="488" reactiontime="+94" swimtime="00:00:28.27" resultid="1292" heatid="3023" lane="8" entrytime="00:00:27.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02016" nation="POL" region="16" clubid="1310" name="Koszalińskie TKKF">
          <ATHLETES>
            <ATHLETE firstname="Marian" lastname="Lasowy" birthdate="1955-07-15" gender="M" nation="POL" license="502016700001" swrid="4967127" athleteid="1322">
              <RESULTS>
                <RESULT eventid="1107" points="115" reactiontime="+103" swimtime="00:03:29.71" resultid="1323" heatid="2998" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                    <SPLIT distance="100" swimtime="00:01:42.90" />
                    <SPLIT distance="150" swimtime="00:02:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="116" reactiontime="+109" swimtime="00:07:30.94" resultid="1324" heatid="3076" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.07" />
                    <SPLIT distance="100" swimtime="00:01:46.60" />
                    <SPLIT distance="150" swimtime="00:02:43.41" />
                    <SPLIT distance="200" swimtime="00:03:41.70" />
                    <SPLIT distance="250" swimtime="00:04:40.11" />
                    <SPLIT distance="300" swimtime="00:05:38.89" />
                    <SPLIT distance="350" swimtime="00:06:36.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lidia" lastname="Mikołajczyk" birthdate="1987-04-29" gender="F" nation="POL" license="102016600013" athleteid="1311">
              <RESULTS>
                <RESULT eventid="1071" points="338" reactiontime="+92" swimtime="00:00:33.96" resultid="1312" heatid="2951" lane="1" />
                <RESULT eventid="1135" points="339" reactiontime="+101" swimtime="00:01:14.14" resultid="1313" heatid="3029" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Mamrot" birthdate="1972-12-10" gender="M" nation="POL" license="102016700007" athleteid="1318">
              <RESULTS>
                <RESULT eventid="1075" points="213" reactiontime="+89" swimtime="00:00:35.01" resultid="1319" heatid="2965" lane="0" />
                <RESULT eventid="1115" points="176" reactiontime="+114" swimtime="00:01:41.40" resultid="1320" heatid="3006" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="198" reactiontime="+94" swimtime="00:00:44.48" resultid="1321" heatid="3052" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Paziewska" birthdate="1974-09-05" gender="F" nation="POL" license="102016600012" athleteid="1314">
              <RESULTS>
                <RESULT eventid="1071" points="317" reactiontime="+86" swimtime="00:00:34.68" resultid="1315" heatid="2954" lane="0" />
                <RESULT eventid="1103" points="272" reactiontime="+100" swimtime="00:02:54.34" resultid="1316" heatid="2996" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:21.68" />
                    <SPLIT distance="150" swimtime="00:02:09.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="308" reactiontime="+92" swimtime="00:01:16.53" resultid="1317" heatid="3029" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01507" nation="POL" region="07" clubid="2631" name="UKS MOS w Opolu">
          <ATHLETES>
            <ATHLETE firstname="Kacper" lastname="Wasztyl" birthdate="2008-04-18" gender="M" nation="POL" license="101507700064" swrid="5041962" athleteid="2632">
              <RESULTS>
                <RESULT eventid="1083" points="384" reactiontime="+75" swimtime="00:02:53.37" resultid="2633" heatid="2974" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:22.01" />
                    <SPLIT distance="150" swimtime="00:02:07.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="354" reactiontime="+82" swimtime="00:01:20.39" resultid="2634" heatid="3006" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="330" reactiontime="+76" swimtime="00:00:37.52" resultid="2635" heatid="3051" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00116" nation="POL" region="16" clubid="2121" name="MKP Szczecin">
          <ATHLETES>
            <ATHLETE firstname="Robert" lastname="Woźnicki" birthdate="1972-03-18" gender="M" nation="POL" license="500116701396" swrid="4302597" athleteid="2135">
              <RESULTS>
                <RESULT eventid="1147" points="173" reactiontime="+91" swimtime="00:00:46.55" resultid="2136" heatid="3053" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Kowalczyk" birthdate="1974-10-02" gender="M" nation="POL" license="500116701197" swrid="4992788" athleteid="2122">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="2123" heatid="2962" lane="8" />
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="2124" heatid="2999" lane="3" />
                <RESULT eventid="1179" status="DNS" swimtime="00:00:00.00" resultid="2125" heatid="3076" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Serbin" birthdate="1966-08-10" gender="F" nation="POL" license="100116601118" swrid="4302596" athleteid="2130">
              <RESULTS>
                <RESULT eventid="1103" points="406" reactiontime="+77" swimtime="00:02:32.49" resultid="2131" heatid="2994" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:13.72" />
                    <SPLIT distance="150" swimtime="00:01:53.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="411" reactiontime="+76" swimtime="00:05:17.95" resultid="2132" heatid="3074" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:16.14" />
                    <SPLIT distance="150" swimtime="00:01:56.35" />
                    <SPLIT distance="200" swimtime="00:02:36.92" />
                    <SPLIT distance="250" swimtime="00:03:17.45" />
                    <SPLIT distance="300" swimtime="00:03:58.16" />
                    <SPLIT distance="350" swimtime="00:04:38.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Szozda" birthdate="1960-01-12" gender="M" nation="POL" license="100116701117" swrid="4461547" athleteid="2126">
              <RESULTS>
                <RESULT eventid="1091" points="150" reactiontime="+134" swimtime="00:01:33.03" resultid="2127" heatid="2981" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="216" reactiontime="+100" swimtime="00:00:37.06" resultid="2128" heatid="3020" lane="5" />
                <RESULT eventid="1147" points="226" reactiontime="+109" swimtime="00:00:42.54" resultid="2129" heatid="3053" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sławomir" lastname="Grzeszewski" birthdate="1953-09-25" gender="M" nation="POL" license="500116701057" swrid="4754656" athleteid="2133">
              <RESULTS>
                <RESULT eventid="1147" points="202" reactiontime="+77" swimtime="00:00:44.18" resultid="2134" heatid="3051" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03914" nation="POL" region="14" clubid="2224" name="Mokotowski UKP Warszawianka- Wodny Park">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Szwedzki" birthdate="2000-12-12" gender="M" nation="POL" license="103914700163" swrid="4001538" athleteid="2225">
              <RESULTS>
                <RESULT eventid="1075" points="496" reactiontime="+75" swimtime="00:00:26.41" resultid="2226" heatid="2962" lane="4" />
                <RESULT eventid="1099" points="426" reactiontime="+74" swimtime="00:00:31.88" resultid="2227" heatid="2990" lane="3" />
                <RESULT eventid="1123" points="432" reactiontime="+71" swimtime="00:00:29.44" resultid="2228" heatid="3022" lane="5" entrytime="00:00:29.25" entrycourse="LCM" />
                <RESULT eventid="1147" points="497" reactiontime="+83" swimtime="00:00:32.76" resultid="2229" heatid="3054" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03715" nation="POL" region="15" clubid="1187" name="&apos;&apos;UKS - Jedynka Kórnik&apos;&apos;">
          <ATHLETES>
            <ATHLETE firstname="Zuzanna" lastname="Deneka" birthdate="2009-01-26" gender="F" nation="POL" license="103715600022" swrid="5334901" athleteid="1202">
              <RESULTS>
                <RESULT eventid="1111" points="283" reactiontime="+70" swimtime="00:01:37.58" resultid="1203" heatid="3004" lane="9" entrytime="00:01:36.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="301" reactiontime="+76" swimtime="00:00:43.83" resultid="1204" heatid="3047" lane="3" entrytime="00:00:44.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nataniel" lastname="Kanikowski" birthdate="2011-10-07" gender="M" nation="POL" license="103715700033" swrid="5448935" athleteid="1192">
              <RESULTS>
                <RESULT eventid="1075" points="169" reactiontime="+60" swimtime="00:00:37.80" resultid="1193" heatid="2965" lane="6" entrytime="00:00:38.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Borys" lastname="Adamczyk" birthdate="2008-04-09" gender="M" nation="POL" license="103715700030" swrid="5448027" athleteid="1190">
              <RESULTS>
                <RESULT eventid="1075" points="367" swimtime="00:00:29.18" resultid="1191" heatid="2967" lane="2" entrytime="00:00:29.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Mocny" birthdate="2010-08-16" gender="M" nation="POL" license="103715700031" swrid="5448037" athleteid="1205">
              <RESULTS>
                <RESULT eventid="1115" points="201" swimtime="00:01:37.07" resultid="1206" heatid="3008" lane="1" entrytime="00:01:34.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="206" reactiontime="+73" swimtime="00:00:43.92" resultid="1207" heatid="3055" lane="1" entrytime="00:00:43.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ignacy" lastname="Rogacki" birthdate="2007-01-15" gender="M" nation="POL" license="103715700026" swrid="5448194" athleteid="1208">
              <RESULTS>
                <RESULT eventid="1147" points="257" swimtime="00:00:40.79" resultid="1209" heatid="3052" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Jabłońska" birthdate="2007-05-10" gender="F" nation="POL" license="103715600014" swrid="5356132" athleteid="1188">
              <RESULTS>
                <RESULT eventid="1071" points="309" reactiontime="+69" swimtime="00:00:35.00" resultid="1189" heatid="2953" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Rogacki" birthdate="2007-07-30" gender="M" nation="POL" license="103715700024" swrid="5443307" athleteid="1194">
              <RESULTS>
                <RESULT eventid="1075" points="260" reactiontime="+51" swimtime="00:00:32.75" resultid="1195" heatid="2960" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Kolba" birthdate="2008-12-09" gender="M" nation="POL" license="103715700032" swrid="5334910" athleteid="1199">
              <RESULTS>
                <RESULT eventid="1099" points="276" reactiontime="+75" swimtime="00:00:36.85" resultid="1200" heatid="2991" lane="7" entrytime="00:00:36.82" entrycourse="LCM" />
                <RESULT eventid="1163" points="282" reactiontime="+85" swimtime="00:01:19.03" resultid="1201" heatid="3064" lane="2" entrytime="00:01:19.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kułton" birthdate="2007-10-09" gender="M" nation="POL" license="103715700011" swrid="5249563" athleteid="1196">
              <RESULTS>
                <RESULT eventid="1091" points="363" reactiontime="+74" swimtime="00:01:09.34" resultid="1197" heatid="2981" lane="6" entrytime="00:01:09.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="409" swimtime="00:00:30.00" resultid="1198" heatid="3022" lane="2" entrytime="00:00:30.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02602" nation="POL" region="02" clubid="2405" name="Toruń Multisport Team">
          <ATHLETES>
            <ATHLETE firstname="Arkadiusz" lastname="Doliński" birthdate="1978-02-06" gender="M" nation="POL" license="502602700088" swrid="4992677" athleteid="2406">
              <RESULTS>
                <RESULT eventid="1075" points="322" reactiontime="+99" swimtime="00:00:30.49" resultid="2407" heatid="2962" lane="9" />
                <RESULT eventid="1099" points="297" reactiontime="+79" swimtime="00:00:35.97" resultid="2408" heatid="2990" lane="6" />
                <RESULT eventid="1123" points="233" reactiontime="+96" swimtime="00:00:36.15" resultid="2409" heatid="3020" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00202" nation="POL" region="02" clubid="2188" name="MKS SP 63 Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Aleksander" lastname="Daniel" birthdate="2007-10-02" gender="M" nation="POL" license="100202700210" swrid="5087014" athleteid="2218">
              <RESULTS>
                <RESULT eventid="1123" points="228" reactiontime="+68" swimtime="00:00:36.45" resultid="2219" heatid="3020" lane="4" />
                <RESULT eventid="1139" points="267" swimtime="00:01:12.76" resultid="2220" heatid="3038" lane="2" entrytime="00:01:13.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Lewicki" birthdate="2007-07-31" gender="M" nation="POL" license="100202700221" swrid="5255261" athleteid="2196">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="2197" heatid="2960" lane="2" />
                <RESULT eventid="1123" points="151" reactiontime="+96" swimtime="00:00:41.76" resultid="2198" heatid="3017" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michalina" lastname="Woźniak" birthdate="2007-08-08" gender="F" nation="POL" license="100202600212" swrid="5087008" athleteid="2207">
              <RESULTS>
                <RESULT eventid="1119" points="483" reactiontime="+73" swimtime="00:00:31.13" resultid="2209" heatid="3012" lane="0" />
                <RESULT eventid="1143" points="501" reactiontime="+82" swimtime="00:00:37.01" resultid="2210" heatid="3045" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Fojutowski" birthdate="2008-10-07" gender="M" nation="POL" license="100202700230" swrid="5163950" athleteid="2221">
              <RESULTS>
                <RESULT eventid="1123" points="312" reactiontime="+61" swimtime="00:00:32.81" resultid="2222" heatid="3018" lane="3" />
                <RESULT eventid="1131" points="261" reactiontime="+61" swimtime="00:02:55.03" resultid="2223" heatid="3027" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:26.27" />
                    <SPLIT distance="150" swimtime="00:02:12.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Rydyńska" birthdate="2007-03-23" gender="F" nation="POL" license="100202600196" swrid="4936885" athleteid="2211">
              <RESULTS>
                <RESULT eventid="1095" points="477" reactiontime="+99" swimtime="00:00:34.53" resultid="2212" heatid="2985" lane="9" />
                <RESULT eventid="1119" points="404" reactiontime="+85" swimtime="00:00:33.04" resultid="2213" heatid="3011" lane="5" />
                <RESULT eventid="1167" points="449" reactiontime="+85" swimtime="00:02:44.69" resultid="2214" heatid="3066" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:01:18.18" />
                    <SPLIT distance="150" swimtime="00:02:08.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sonia" lastname="Matuszyńska" birthdate="2006-06-19" gender="F" nation="POL" license="100202600185" swrid="4933946" athleteid="2189">
              <RESULTS>
                <RESULT eventid="1071" points="478" reactiontime="+72" swimtime="00:00:30.27" resultid="2190" heatid="2957" lane="1" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1135" points="462" reactiontime="+69" swimtime="00:01:06.86" resultid="2191" heatid="3032" lane="5" entrytime="00:01:06.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="437" reactiontime="+74" swimtime="00:02:46.09" resultid="2192" heatid="3066" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:18.57" />
                    <SPLIT distance="150" swimtime="00:02:08.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Franciszek" lastname="Bakalarz" birthdate="2007-09-16" gender="M" nation="POL" license="100202700211" swrid="5087013" athleteid="2193">
              <RESULTS>
                <RESULT eventid="1075" points="406" reactiontime="+72" swimtime="00:00:28.23" resultid="2194" heatid="2968" lane="6" entrytime="00:00:27.90" entrycourse="LCM" />
                <RESULT eventid="1123" points="403" reactiontime="+75" swimtime="00:00:30.13" resultid="2195" heatid="3020" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Fojutowski" birthdate="2006-03-22" gender="M" nation="POL" license="100202700145" swrid="4997751" athleteid="2199">
              <RESULTS>
                <RESULT eventid="1075" points="372" reactiontime="+64" swimtime="00:00:29.05" resultid="2200" heatid="2968" lane="1" entrytime="00:00:28.49" entrycourse="LCM" />
                <RESULT eventid="1123" points="290" reactiontime="+69" swimtime="00:00:33.61" resultid="2201" heatid="3020" lane="8" />
                <RESULT eventid="1147" points="292" reactiontime="+76" swimtime="00:00:39.10" resultid="2202" heatid="3054" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Ławrynowicz" birthdate="2009-07-14" gender="M" nation="POL" license="100202700243" swrid="5042257" athleteid="2203">
              <RESULTS>
                <RESULT eventid="1083" points="257" swimtime="00:03:18.14" resultid="2204" heatid="2974" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                    <SPLIT distance="100" swimtime="00:01:34.31" />
                    <SPLIT distance="150" swimtime="00:02:26.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="277" reactiontime="+61" swimtime="00:00:34.15" resultid="2205" heatid="3021" lane="9" />
                <RESULT eventid="1171" points="279" reactiontime="+77" swimtime="00:02:54.34" resultid="2206" heatid="3070" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:01:24.19" />
                    <SPLIT distance="150" swimtime="00:02:15.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Ratajczak" birthdate="2008-05-20" gender="M" nation="POL" license="100202700232" swrid="5108575" athleteid="2215">
              <RESULTS>
                <RESULT eventid="1099" points="297" reactiontime="+61" swimtime="00:00:35.97" resultid="2216" heatid="2991" lane="6" entrytime="00:00:35.70" entrycourse="LCM" />
                <RESULT eventid="1131" points="271" reactiontime="+67" swimtime="00:02:52.88" resultid="2217" heatid="3028" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:26.19" />
                    <SPLIT distance="150" swimtime="00:02:12.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03102" nation="POL" region="02" clubid="2382" name="St. KP Olimpia Świecie">
          <ATHLETES>
            <ATHLETE firstname="Alicja" lastname="Szczepańska" birthdate="2005-11-09" gender="F" nation="POL" license="103102600033" swrid="4924065" athleteid="2388">
              <RESULTS>
                <RESULT eventid="1071" points="565" reactiontime="+63" swimtime="00:00:28.63" resultid="2389" heatid="2959" lane="1" entrytime="00:00:28.19" entrycourse="LCM" />
                <RESULT eventid="1087" points="478" reactiontime="+62" swimtime="00:01:10.92" resultid="2390" heatid="2979" lane="0" entrytime="00:01:08.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="507" reactiontime="+74" swimtime="00:00:33.82" resultid="2391" heatid="2986" lane="4" entrytime="00:00:35.13" entrycourse="LCM" />
                <RESULT eventid="1119" points="491" reactiontime="+63" swimtime="00:00:30.95" resultid="2392" heatid="3015" lane="3" entrytime="00:00:31.10" entrycourse="LCM" />
                <RESULT eventid="1135" points="540" reactiontime="+62" swimtime="00:01:03.49" resultid="2393" heatid="3034" lane="0" entrytime="00:01:01.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Klonowski" birthdate="2007-12-19" gender="M" nation="POL" license="103102700006" swrid="4923763" athleteid="2383">
              <RESULTS>
                <RESULT eventid="1099" points="349" reactiontime="+64" swimtime="00:00:34.07" resultid="2385" heatid="2988" lane="6" />
                <RESULT eventid="1131" points="395" reactiontime="+60" swimtime="00:02:32.45" resultid="2386" heatid="3028" lane="2" entrytime="00:02:33.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:14.79" />
                    <SPLIT distance="150" swimtime="00:01:54.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="375" reactiontime="+62" swimtime="00:01:11.85" resultid="2387" heatid="3064" lane="4" entrytime="00:01:12.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1091" points="265" reactiontime="+69" swimtime="00:01:17.05" resultid="2810" heatid="2980" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Hofman" birthdate="2008-03-14" gender="M" nation="POL" license="100802700370" swrid="4923739" athleteid="2394">
              <RESULTS>
                <RESULT eventid="1075" points="292" reactiontime="+75" swimtime="00:00:31.50" resultid="2395" heatid="2966" lane="3" entrytime="00:00:30.92" entrycourse="LCM" />
                <RESULT eventid="1099" points="239" reactiontime="+75" swimtime="00:00:38.62" resultid="2396" heatid="2991" lane="0" entrytime="00:00:39.09" entrycourse="LCM" />
                <RESULT eventid="1123" points="225" reactiontime="+82" swimtime="00:00:36.57" resultid="2397" heatid="3019" lane="7" />
                <RESULT eventid="1147" points="178" reactiontime="+76" swimtime="00:00:46.09" resultid="2398" heatid="3053" lane="8" />
                <RESULT eventid="1171" points="236" reactiontime="+81" swimtime="00:03:04.40" resultid="2399" heatid="3071" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.20" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                    <SPLIT distance="150" swimtime="00:02:24.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03302" nation="POL" region="02" clubid="2410" name="Toruński MKS CHAMPIONS">
          <ATHLETES>
            <ATHLETE firstname="Kazimierz" lastname="Piotrowski" birthdate="1952-12-22" gender="M" nation="POL" license="103302700073" swrid="5337365" athleteid="2411">
              <RESULTS>
                <RESULT eventid="1075" points="103" reactiontime="+107" swimtime="00:00:44.47" resultid="2412" heatid="2965" lane="7" entrytime="00:00:43.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02101" nation="POL" region="01" clubid="2426" name="UKS &apos;&apos;ORKA&apos;&apos; Lubań">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Kozik" birthdate="2006-04-19" gender="M" nation="POL" license="102101700060" swrid="5024309" athleteid="2435">
              <RESULTS>
                <RESULT eventid="1075" points="547" reactiontime="+74" swimtime="00:00:25.56" resultid="2436" heatid="2970" lane="4" entrytime="00:00:25.42" entrycourse="LCM" />
                <RESULT eventid="1123" points="502" swimtime="00:00:28.02" resultid="2437" heatid="3023" lane="2" entrytime="00:00:27.62" entrycourse="LCM" />
                <RESULT eventid="1139" points="541" reactiontime="+71" swimtime="00:00:57.57" resultid="2438" heatid="3042" lane="6" entrytime="00:00:56.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Wasyliszyn" birthdate="2004-04-26" gender="F" nation="POL" license="102101600062" swrid="5094195" athleteid="2427">
              <RESULTS>
                <RESULT eventid="1071" points="403" reactiontime="+78" swimtime="00:00:32.02" resultid="2428" heatid="2951" lane="0" />
                <RESULT eventid="1111" points="378" reactiontime="+89" swimtime="00:01:28.67" resultid="2429" heatid="3002" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="381" reactiontime="+82" swimtime="00:00:40.52" resultid="2430" heatid="3045" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julita" lastname="Jośko" birthdate="2004-04-30" gender="F" nation="POL" license="102101600129" swrid="4910964" athleteid="2431">
              <RESULTS>
                <RESULT eventid="1071" points="506" reactiontime="+69" swimtime="00:00:29.69" resultid="2432" heatid="2957" lane="0" entrytime="00:00:30.05" entrycourse="LCM" />
                <RESULT eventid="1095" points="463" reactiontime="+79" swimtime="00:00:34.85" resultid="2433" heatid="2986" lane="3" entrytime="00:00:35.19" entrycourse="LCM" />
                <RESULT eventid="1159" points="402" reactiontime="+77" swimtime="00:01:17.96" resultid="2434" heatid="3061" lane="3" entrytime="00:01:17.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02815" nation="POL" region="15" clubid="2439" name="UKS ,,GROT&apos;&apos; Koziegłowy">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Mizerska" birthdate="2006-06-16" gender="F" nation="POL" license="102815600104" swrid="4975736" athleteid="2440">
              <RESULTS>
                <RESULT eventid="1119" points="228" reactiontime="+88" swimtime="00:00:39.97" resultid="2441" heatid="3012" lane="3" />
                <RESULT eventid="1143" points="297" reactiontime="+75" swimtime="00:00:44.06" resultid="2442" heatid="3045" lane="5" />
                <RESULT eventid="1167" points="299" reactiontime="+87" swimtime="00:03:08.40" resultid="2443" heatid="3067" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:31.18" />
                    <SPLIT distance="150" swimtime="00:02:25.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02305" nation="POL" region="05" clubid="1257" name="AZS UŁ PŁ Łódź">
          <ATHLETES>
            <ATHLETE firstname="Wiktoria" lastname="Raczyńska" birthdate="2004-04-16" gender="F" nation="POL" license="102305600064" swrid="5034876" athleteid="1258">
              <RESULTS>
                <RESULT eventid="1071" points="494" swimtime="00:00:29.93" resultid="1259" heatid="2957" lane="2" entrytime="00:00:29.76" entrycourse="LCM" />
                <RESULT eventid="1087" points="542" reactiontime="+70" swimtime="00:01:08.01" resultid="1260" heatid="2979" lane="1" entrytime="00:01:07.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="486" reactiontime="+70" swimtime="00:00:31.06" resultid="1261" heatid="3016" lane="7" entrytime="00:00:29.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06115" nation="POL" region="15" clubid="1210" name="Aquapark Wągrowiec sp. z o.o.">
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Spychalska" birthdate="2008-06-06" gender="F" nation="POL" license="106115600025" swrid="4865406" athleteid="1239">
              <RESULTS>
                <RESULT eventid="1103" points="351" reactiontime="+108" swimtime="00:02:40.15" resultid="1240" heatid="2996" lane="7" entrytime="00:02:31.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="150" swimtime="00:02:00.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="326" reactiontime="+98" swimtime="00:02:59.19" resultid="1241" heatid="3026" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                    <SPLIT distance="100" swimtime="00:01:30.07" />
                    <SPLIT distance="150" swimtime="00:02:16.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="331" reactiontime="+91" swimtime="00:05:41.67" resultid="1242" heatid="3074" lane="7" entrytime="00:05:25.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:01:21.39" />
                    <SPLIT distance="150" swimtime="00:02:05.47" />
                    <SPLIT distance="200" swimtime="00:02:49.16" />
                    <SPLIT distance="250" swimtime="00:03:33.31" />
                    <SPLIT distance="300" swimtime="00:04:17.80" />
                    <SPLIT distance="350" swimtime="00:05:01.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Pilarska" birthdate="2008-12-15" gender="F" nation="POL" license="106115600018" swrid="5190193" athleteid="1225">
              <RESULTS>
                <RESULT eventid="1079" points="301" reactiontime="+86" swimtime="00:03:27.56" resultid="1226" heatid="2972" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                    <SPLIT distance="100" swimtime="00:01:41.19" />
                    <SPLIT distance="150" swimtime="00:02:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="260" swimtime="00:01:40.44" resultid="1227" heatid="3002" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="239" swimtime="00:00:47.31" resultid="1228" heatid="3047" lane="2" entrytime="00:00:45.56" entrycourse="LCM" />
                <RESULT eventid="1167" points="266" reactiontime="+59" swimtime="00:03:16.09" resultid="1229" heatid="3068" lane="9" entrytime="00:03:06.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                    <SPLIT distance="100" swimtime="00:01:36.51" />
                    <SPLIT distance="150" swimtime="00:02:30.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Paszek" birthdate="2008-03-03" gender="M" nation="POL" license="106115700010" swrid="5448915" athleteid="1216">
              <RESULTS>
                <RESULT eventid="1075" points="263" reactiontime="+86" swimtime="00:00:32.60" resultid="1217" heatid="2966" lane="1" entrytime="00:00:32.04" entrycourse="LCM" />
                <RESULT eventid="1099" points="213" reactiontime="+88" swimtime="00:00:40.18" resultid="1218" heatid="2991" lane="9" entrytime="00:00:39.68" entrycourse="LCM" />
                <RESULT eventid="1107" points="260" reactiontime="+80" swimtime="00:02:39.70" resultid="1219" heatid="3000" lane="0" entrytime="00:02:42.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="150" swimtime="00:01:57.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="265" reactiontime="+65" swimtime="00:01:12.97" resultid="1220" heatid="3038" lane="5" entrytime="00:01:11.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Starzyński" birthdate="2006-04-20" gender="M" nation="POL" license="106115700014" swrid="5190202" athleteid="1235">
              <RESULTS>
                <RESULT eventid="1099" points="519" reactiontime="+59" swimtime="00:00:29.86" resultid="1236" heatid="2992" lane="5" entrytime="00:00:29.84" entrycourse="LCM" />
                <RESULT eventid="1131" points="444" reactiontime="+61" swimtime="00:02:26.64" resultid="1237" heatid="3028" lane="7" entrytime="00:02:39.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:09.70" />
                    <SPLIT distance="150" swimtime="00:01:47.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="492" reactiontime="+58" swimtime="00:01:05.64" resultid="1238" heatid="3065" lane="0" entrytime="00:01:06.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Chomko" birthdate="2008-08-11" gender="F" nation="POL" license="106115600021" swrid="4722169" athleteid="1211">
              <RESULTS>
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="1212" heatid="2953" lane="6" />
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="1213" heatid="2972" lane="1" />
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="1214" heatid="3004" lane="8" entrytime="00:01:32.77" entrycourse="LCM" />
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="1215" heatid="3048" lane="9" entrytime="00:00:43.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Makarewicz" birthdate="2006-06-16" gender="M" nation="POL" license="106115700012" swrid="4865304" athleteid="1243">
              <RESULTS>
                <RESULT eventid="1107" points="491" reactiontime="+65" swimtime="00:02:09.28" resultid="1244" heatid="3001" lane="1" entrytime="00:02:09.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:02.43" />
                    <SPLIT distance="150" swimtime="00:01:36.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="454" reactiontime="+67" swimtime="00:04:46.15" resultid="1245" heatid="3077" lane="3" entrytime="00:04:41.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:07.56" />
                    <SPLIT distance="150" swimtime="00:01:44.80" />
                    <SPLIT distance="200" swimtime="00:02:22.41" />
                    <SPLIT distance="250" swimtime="00:02:59.24" />
                    <SPLIT distance="300" swimtime="00:03:36.69" />
                    <SPLIT distance="350" swimtime="00:04:12.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Franciszek" lastname="Drewicz" birthdate="2009-07-18" gender="M" nation="POL" license="106115700109" swrid="5340956" athleteid="1221">
              <RESULTS>
                <RESULT eventid="1075" points="135" reactiontime="+94" swimtime="00:00:40.73" resultid="1222" heatid="2963" lane="8" />
                <RESULT eventid="1099" points="109" reactiontime="+83" swimtime="00:00:50.17" resultid="1223" heatid="2989" lane="2" />
                <RESULT eventid="1147" points="116" reactiontime="+78" swimtime="00:00:53.17" resultid="1224" heatid="3053" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Łatka" birthdate="2008-10-15" gender="M" nation="POL" license="106115700026" swrid="5190194" athleteid="1246">
              <RESULTS>
                <RESULT eventid="1107" points="214" swimtime="00:02:50.50" resultid="1247" heatid="2999" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:22.11" />
                    <SPLIT distance="150" swimtime="00:02:06.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="176" swimtime="00:01:41.39" resultid="1248" heatid="3006" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="164" reactiontime="+78" swimtime="00:00:47.34" resultid="1249" heatid="3051" lane="6" />
                <RESULT eventid="1179" points="198" reactiontime="+96" swimtime="00:06:17.06" resultid="1250" heatid="3076" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                    <SPLIT distance="100" swimtime="00:01:30.49" />
                    <SPLIT distance="150" swimtime="00:02:18.64" />
                    <SPLIT distance="200" swimtime="00:03:06.83" />
                    <SPLIT distance="250" swimtime="00:03:55.76" />
                    <SPLIT distance="300" swimtime="00:04:44.09" />
                    <SPLIT distance="350" swimtime="00:05:32.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1059" swimtime="00:02:15.85" resultid="1251" heatid="2948" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="100" swimtime="00:01:07.82" />
                    <SPLIT distance="150" swimtime="00:01:43.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1216" number="1" />
                    <RELAYPOSITION athleteid="1225" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="1246" number="3" />
                    <RELAYPOSITION athleteid="1239" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="11" clubid="2374" name="AZS AWF Katowice">
          <ATHLETES>
            <ATHLETE firstname="Matylda" lastname="Tuszyńska" birthdate="2005-10-17" gender="F" nation="POL" license="100611600365" swrid="5116172" athleteid="2375">
              <RESULTS>
                <RESULT eventid="1071" points="495" reactiontime="+78" swimtime="00:00:29.91" resultid="2376" heatid="2957" lane="6" entrytime="00:00:29.56" entrycourse="LCM" />
                <RESULT eventid="1159" points="538" reactiontime="+83" swimtime="00:01:10.75" resultid="2377" heatid="3062" lane="8" entrytime="00:01:10.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iga" lastname="Idzikowska" birthdate="2005-04-03" gender="F" nation="POL" license="100611600362" swrid="5057160" athleteid="2378">
              <RESULTS>
                <RESULT eventid="1079" points="584" reactiontime="+65" swimtime="00:02:46.36" resultid="2379" heatid="2973" lane="5" entrytime="00:02:43.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                    <SPLIT distance="100" swimtime="00:01:22.57" />
                    <SPLIT distance="150" swimtime="00:02:05.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="554" reactiontime="+84" swimtime="00:01:18.05" resultid="2380" heatid="3005" lane="3" entrytime="00:01:15.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="506" reactiontime="+87" swimtime="00:02:38.18" resultid="2381" heatid="3067" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                    <SPLIT distance="100" swimtime="00:01:16.65" />
                    <SPLIT distance="150" swimtime="00:02:00.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02805" nation="POL" region="05" clubid="2363" name="MUKS Zgierz">
          <ATHLETES>
            <ATHLETE firstname="Grzegorz" lastname="Januszkiewicz" birthdate="1959-02-19" gender="M" nation="POL" license="502805700130" athleteid="2364">
              <RESULTS>
                <RESULT eventid="1075" points="182" reactiontime="+118" swimtime="00:00:36.85" resultid="2365" heatid="2964" lane="0" />
                <RESULT eventid="1099" points="149" reactiontime="+86" swimtime="00:00:45.25" resultid="2366" heatid="2988" lane="5" />
                <RESULT eventid="1123" points="116" reactiontime="+105" swimtime="00:00:45.58" resultid="2367" heatid="3018" lane="5" />
                <RESULT eventid="1139" points="153" reactiontime="+116" swimtime="00:01:27.65" resultid="2368" heatid="3037" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08114" nation="POL" region="14" clubid="1253" name="AZS  KU Uniwersytetu Warszawskiego">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Micorek" birthdate="1993-08-25" gender="M" nation="POL" license="108114700041" swrid="4086676" athleteid="1254">
              <RESULTS>
                <RESULT eventid="1091" points="479" reactiontime="+91" swimtime="00:01:03.25" resultid="1255" heatid="2980" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02201" nation="POL" region="01" clubid="2662" name="UKS Shark Rudna">
          <ATHLETES>
            <ATHLETE firstname="Szymon" lastname="Misiak" birthdate="2005-12-14" gender="M" nation="POL" license="102201700081" swrid="5135289" athleteid="2668">
              <RESULTS>
                <RESULT eventid="1075" points="633" reactiontime="+73" swimtime="00:00:24.35" resultid="2669" heatid="2971" lane="3" entrytime="00:00:24.11" entrycourse="LCM" />
                <RESULT eventid="1091" points="564" reactiontime="+68" swimtime="00:00:59.88" resultid="2670" heatid="2982" lane="5" entrytime="00:00:58.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="624" reactiontime="+72" swimtime="00:00:26.06" resultid="2671" heatid="3024" lane="6" entrytime="00:00:25.61" entrycourse="LCM" />
                <RESULT eventid="1139" points="622" reactiontime="+73" swimtime="00:00:54.94" resultid="2672" heatid="3043" lane="4" entrytime="00:00:54.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Trzpil" birthdate="2005-03-17" gender="M" nation="POL" license="102201700084" swrid="5148198" athleteid="2673">
              <RESULTS>
                <RESULT eventid="1075" points="537" reactiontime="+73" swimtime="00:00:25.71" resultid="2674" heatid="2970" lane="6" entrytime="00:00:25.58" entrycourse="LCM" />
                <RESULT eventid="1091" points="496" reactiontime="+77" swimtime="00:01:02.52" resultid="2675" heatid="2980" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="452" reactiontime="+80" swimtime="00:01:14.09" resultid="2676" heatid="3009" lane="3" entrytime="00:01:11.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="455" reactiontime="+73" swimtime="00:00:33.73" resultid="2677" heatid="3056" lane="4" entrytime="00:00:32.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Kościelniak" birthdate="2002-06-07" gender="F" nation="POL" license="102201600063" swrid="4892800" athleteid="2663">
              <RESULTS>
                <RESULT eventid="1071" points="606" reactiontime="+74" swimtime="00:00:27.97" resultid="2664" heatid="2959" lane="7" entrytime="00:00:27.93" entrycourse="LCM" />
                <RESULT eventid="1087" points="613" reactiontime="+78" swimtime="00:01:05.30" resultid="2665" heatid="2979" lane="4" entrytime="00:01:05.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="637" reactiontime="+67" swimtime="00:00:28.38" resultid="2666" heatid="3016" lane="5" entrytime="00:00:28.12" entrycourse="LCM" />
                <RESULT eventid="1159" points="629" reactiontime="+52" swimtime="00:01:07.17" resultid="2667" heatid="3062" lane="5" entrytime="00:01:07.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Adamczewska" birthdate="2004-04-06" gender="F" nation="POL" license="102201600092" swrid="5024285" athleteid="2678">
              <RESULTS>
                <RESULT eventid="1087" points="552" reactiontime="+71" swimtime="00:01:07.61" resultid="2679" heatid="2978" lane="4" entrytime="00:01:08.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="533" reactiontime="+43" swimtime="00:01:19.07" resultid="2680" heatid="3005" lane="2" entrytime="00:01:18.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="551" reactiontime="+73" swimtime="00:00:35.85" resultid="2681" heatid="3049" lane="7" entrytime="00:00:35.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adela" lastname="Piskorska" birthdate="2003-11-16" gender="F" nation="POL" license="102201600099" swrid="4931147" athleteid="2682">
              <RESULTS>
                <RESULT eventid="1095" points="806" reactiontime="+61" swimtime="00:00:28.98" resultid="2683" heatid="2987" lane="4" entrytime="00:00:28.78" entrycourse="LCM" />
                <RESULT eventid="1159" points="789" reactiontime="+61" swimtime="00:01:02.28" resultid="2684" heatid="3062" lane="4" entrytime="00:01:01.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="661" reactiontime="+70" swimtime="00:02:24.75" resultid="2685" heatid="3068" lane="5" entrytime="00:02:32.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                    <SPLIT distance="150" swimtime="00:01:51.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04915" nation="POL" region="15" clubid="1301" name="Klub Sportowy Extreme Team Oborniki">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Wolniewicz" birthdate="1948-12-22" gender="M" nation="POL" license="504915700022" swrid="4754624" athleteid="1302">
              <RESULTS>
                <RESULT eventid="1107" points="97" reactiontime="+112" swimtime="00:03:41.81" resultid="1303" heatid="2999" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.87" />
                    <SPLIT distance="100" swimtime="00:01:39.97" />
                    <SPLIT distance="150" swimtime="00:02:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="90" reactiontime="+81" swimtime="00:08:10.94" resultid="1304" heatid="3075" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.79" />
                    <SPLIT distance="100" swimtime="00:01:53.78" />
                    <SPLIT distance="150" swimtime="00:02:56.05" />
                    <SPLIT distance="200" swimtime="00:04:01.16" />
                    <SPLIT distance="250" swimtime="00:05:05.72" />
                    <SPLIT distance="300" swimtime="00:06:10.22" />
                    <SPLIT distance="350" swimtime="00:07:11.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01102" nation="POL" region="02" clubid="2650" name="UKS Ruch Grudziądz">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Zawadzki" birthdate="2006-05-16" gender="M" nation="POL" license="101102700014" swrid="5108583" athleteid="2656">
              <RESULTS>
                <RESULT eventid="1099" points="384" reactiontime="+82" swimtime="00:00:33.00" resultid="2657" heatid="2992" lane="9" entrytime="00:00:33.54" entrycourse="LCM" />
                <RESULT eventid="1139" points="425" swimtime="00:01:02.35" resultid="2658" heatid="3039" lane="2" entrytime="00:01:04.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="330" reactiontime="+66" swimtime="00:00:37.55" resultid="2659" heatid="3052" lane="1" />
                <RESULT eventid="1163" points="373" reactiontime="+74" swimtime="00:01:11.99" resultid="2660" heatid="3065" lane="9" entrytime="00:01:11.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="395" reactiontime="+75" swimtime="00:02:35.34" resultid="2661" heatid="3071" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                    <SPLIT distance="150" swimtime="00:01:59.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Malinowska" birthdate="2008-03-21" gender="F" nation="POL" license="101102600022" swrid="5159067" athleteid="2651">
              <RESULTS>
                <RESULT eventid="1079" points="371" reactiontime="+67" swimtime="00:03:13.46" resultid="2652" heatid="2973" lane="1" entrytime="00:03:06.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:01:31.04" />
                    <SPLIT distance="150" swimtime="00:02:21.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="386" reactiontime="+65" swimtime="00:02:35.10" resultid="2653" heatid="2996" lane="8" entrytime="00:02:34.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="150" swimtime="00:01:54.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="401" reactiontime="+60" swimtime="00:01:10.08" resultid="2654" heatid="3032" lane="9" entrytime="00:01:08.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="400" reactiontime="+58" swimtime="00:00:39.90" resultid="2655" heatid="3048" lane="6" entrytime="00:00:39.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01115" nation="POL" region="15" clubid="1305" name="Klub Sportowy Krotosz Krotoszyn">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Bielawna" birthdate="2004-05-23" gender="F" nation="POL" license="101115600066" swrid="4853998" athleteid="1306">
              <RESULTS>
                <RESULT eventid="1079" points="431" reactiontime="+80" swimtime="00:03:04.16" resultid="1307" heatid="2972" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                    <SPLIT distance="100" swimtime="00:01:28.14" />
                    <SPLIT distance="150" swimtime="00:02:17.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="504" reactiontime="+67" swimtime="00:01:20.56" resultid="1308" heatid="3005" lane="0" entrytime="00:01:23.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="536" reactiontime="+73" swimtime="00:00:36.19" resultid="1309" heatid="3049" lane="8" entrytime="00:00:36.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04901" nation="POL" region="01" clubid="1388" name="KS Neptun Świdnica">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Jackowski" birthdate="2002-06-10" gender="M" nation="POL" license="104901700069" swrid="4929919" athleteid="1414">
              <RESULTS>
                <RESULT eventid="1075" points="575" reactiontime="+72" swimtime="00:00:25.14" resultid="1415" heatid="2960" lane="4" />
                <RESULT eventid="1091" points="592" reactiontime="+70" swimtime="00:00:58.92" resultid="1416" heatid="2982" lane="7" entrytime="00:01:01.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="557" reactiontime="+70" swimtime="00:00:27.06" resultid="1417" heatid="3023" lane="7" entrytime="00:00:27.69" entrycourse="LCM" />
                <RESULT eventid="1139" points="662" swimtime="00:00:53.81" resultid="1418" heatid="3043" lane="2" entrytime="00:00:55.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Wrona" birthdate="2008-09-03" gender="F" nation="POL" license="104901600034" swrid="5272089" athleteid="1401">
              <RESULTS>
                <RESULT eventid="1071" points="280" swimtime="00:00:36.18" resultid="1402" heatid="2954" lane="2" entrytime="00:00:36.14" entrycourse="LCM" />
                <RESULT eventid="1111" points="209" swimtime="00:01:48.00" resultid="1403" heatid="3003" lane="5" entrytime="00:01:51.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="198" swimtime="00:00:50.39" resultid="1404" heatid="3047" lane="7" entrytime="00:00:49.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ignacy" lastname="Stachyra" birthdate="2009-09-08" gender="M" nation="POL" license="104901700048" swrid="5395485" athleteid="1434">
              <RESULTS>
                <RESULT eventid="1083" points="230" reactiontime="+87" swimtime="00:03:25.57" resultid="1435" heatid="2974" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.57" />
                    <SPLIT distance="100" swimtime="00:01:40.43" />
                    <SPLIT distance="150" swimtime="00:02:33.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="197" swimtime="00:01:37.70" resultid="1436" heatid="3008" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="210" reactiontime="+85" swimtime="00:00:43.59" resultid="1437" heatid="3055" lane="8" entrytime="00:00:45.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Kuśnierz" birthdate="2006-02-11" gender="F" nation="POL" license="104901600029" swrid="5165939" athleteid="1422">
              <RESULTS>
                <RESULT eventid="1079" points="425" reactiontime="+81" swimtime="00:03:04.99" resultid="1423" heatid="2973" lane="7" entrytime="00:03:05.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                    <SPLIT distance="100" swimtime="00:01:29.16" />
                    <SPLIT distance="150" swimtime="00:02:17.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="408" reactiontime="+88" swimtime="00:01:26.42" resultid="1424" heatid="3005" lane="9" entrytime="00:01:24.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="435" reactiontime="+69" swimtime="00:00:38.80" resultid="1425" heatid="3048" lane="5" entrytime="00:00:37.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Lęga" birthdate="2005-04-20" gender="F" nation="POL" license="104901600009" swrid="4995402" athleteid="1389">
              <RESULTS>
                <RESULT eventid="1071" points="487" reactiontime="+78" swimtime="00:00:30.08" resultid="1390" heatid="2957" lane="5" entrytime="00:00:29.47" entrycourse="LCM" />
                <RESULT eventid="1135" points="498" reactiontime="+72" swimtime="00:01:05.21" resultid="1391" heatid="3033" lane="3" entrytime="00:01:03.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="495" reactiontime="+76" swimtime="00:04:58.92" resultid="1392" heatid="3074" lane="3" entrytime="00:04:56.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:10.73" />
                    <SPLIT distance="150" swimtime="00:01:48.65" />
                    <SPLIT distance="200" swimtime="00:02:26.55" />
                    <SPLIT distance="250" swimtime="00:03:05.10" />
                    <SPLIT distance="300" swimtime="00:03:43.17" />
                    <SPLIT distance="350" swimtime="00:04:21.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Cichoń" birthdate="2009-07-24" gender="M" nation="POL" license="104901700040" swrid="5341304" athleteid="1410">
              <RESULTS>
                <RESULT eventid="1075" points="242" reactiontime="+75" swimtime="00:00:33.52" resultid="1411" heatid="2961" lane="1" />
                <RESULT eventid="1091" points="184" reactiontime="+75" swimtime="00:01:26.98" resultid="1412" heatid="2980" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="257" reactiontime="+78" swimtime="00:01:13.77" resultid="1413" heatid="3038" lane="7" entrytime="00:01:14.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Skroboń" birthdate="2009-10-16" gender="F" nation="POL" license="104901600049" swrid="5449672" athleteid="1430">
              <RESULTS>
                <RESULT eventid="1079" points="318" reactiontime="+79" swimtime="00:03:23.80" resultid="1431" heatid="2972" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="100" swimtime="00:01:39.30" />
                    <SPLIT distance="150" swimtime="00:02:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="296" reactiontime="+83" swimtime="00:01:36.15" resultid="1432" heatid="3003" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="302" reactiontime="+76" swimtime="00:00:43.79" resultid="1433" heatid="3047" lane="6" entrytime="00:00:45.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Oleksy" birthdate="2009-04-04" gender="F" nation="POL" license="104901600041" swrid="5356111" athleteid="1397">
              <RESULTS>
                <RESULT eventid="1071" points="203" reactiontime="+92" swimtime="00:00:40.24" resultid="1398" heatid="2954" lane="8" entrytime="00:00:40.30" entrycourse="LCM" />
                <RESULT eventid="1095" points="172" reactiontime="+78" swimtime="00:00:48.46" resultid="1399" heatid="2985" lane="3" entrytime="00:00:47.80" entrycourse="LCM" />
                <RESULT eventid="1143" points="173" reactiontime="+84" swimtime="00:00:52.75" resultid="1400" heatid="3047" lane="8" entrytime="00:00:58.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Jaros" birthdate="2009-07-18" gender="F" nation="POL" license="104901600042" swrid="5244068" athleteid="1426">
              <RESULTS>
                <RESULT eventid="1079" points="261" reactiontime="+70" swimtime="00:03:37.45" resultid="1427" heatid="2972" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.96" />
                    <SPLIT distance="100" swimtime="00:01:45.98" />
                    <SPLIT distance="150" swimtime="00:02:42.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="253" reactiontime="+77" swimtime="00:01:41.30" resultid="1428" heatid="3003" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="236" reactiontime="+68" swimtime="00:00:47.51" resultid="1429" heatid="3047" lane="1" entrytime="00:00:52.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamila" lastname="Świdnicka" birthdate="2006-06-07" gender="F" nation="POL" license="104901600068" swrid="4995331" athleteid="1438">
              <RESULTS>
                <RESULT eventid="1103" points="540" reactiontime="+74" swimtime="00:02:18.72" resultid="1439" heatid="2997" lane="8" entrytime="00:02:19.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:06.90" />
                    <SPLIT distance="150" swimtime="00:01:43.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="532" reactiontime="+79" swimtime="00:01:03.80" resultid="1440" heatid="3033" lane="6" entrytime="00:01:03.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="535" reactiontime="+77" swimtime="00:04:51.16" resultid="1441" heatid="3074" lane="6" entrytime="00:04:58.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:47.12" />
                    <SPLIT distance="200" swimtime="00:02:24.53" />
                    <SPLIT distance="250" swimtime="00:03:01.81" />
                    <SPLIT distance="300" swimtime="00:03:39.46" />
                    <SPLIT distance="350" swimtime="00:04:16.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Kowalik" birthdate="2006-06-07" gender="M" nation="POL" license="104901700016" swrid="5165949" athleteid="1405">
              <RESULTS>
                <RESULT eventid="1075" points="359" reactiontime="+69" swimtime="00:00:29.40" resultid="1406" heatid="2967" lane="6" entrytime="00:00:29.57" entrycourse="LCM" />
                <RESULT eventid="1107" points="369" reactiontime="+75" swimtime="00:02:22.08" resultid="1407" heatid="3000" lane="2" entrytime="00:02:19.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:07.21" />
                    <SPLIT distance="150" swimtime="00:01:44.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="377" reactiontime="+82" swimtime="00:01:04.91" resultid="1408" heatid="3040" lane="9" entrytime="00:01:02.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="389" reactiontime="+76" swimtime="00:05:01.42" resultid="1409" heatid="3077" lane="7" entrytime="00:04:54.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="150" swimtime="00:01:48.31" />
                    <SPLIT distance="200" swimtime="00:02:27.28" />
                    <SPLIT distance="250" swimtime="00:03:06.17" />
                    <SPLIT distance="300" swimtime="00:03:45.39" />
                    <SPLIT distance="350" swimtime="00:04:24.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Łazarz" birthdate="2006-06-26" gender="F" nation="POL" license="104901600062" swrid="5450902" athleteid="1393">
              <RESULTS>
                <RESULT eventid="1071" points="222" reactiontime="+94" swimtime="00:00:39.09" resultid="1394" heatid="2952" lane="1" />
                <RESULT eventid="1095" points="200" reactiontime="+85" swimtime="00:00:46.09" resultid="1395" heatid="2984" lane="4" />
                <RESULT eventid="1143" points="214" reactiontime="+74" swimtime="00:00:49.13" resultid="1396" heatid="3045" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kinga" lastname="Kamieniarz" birthdate="2005-04-09" gender="F" nation="POL" license="104901600046" swrid="5166049" athleteid="1419">
              <RESULTS>
                <RESULT eventid="1079" points="617" reactiontime="+67" swimtime="00:02:43.40" resultid="1420" heatid="2973" lane="3" entrytime="00:02:44.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:19.79" />
                    <SPLIT distance="150" swimtime="00:02:01.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="578" reactiontime="+66" swimtime="00:01:16.95" resultid="1421" heatid="3005" lane="6" entrytime="00:01:17.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04115" nation="POL" region="15" clubid="1888" name="KTP Iskra Konin">
          <ATHLETES>
            <ATHLETE firstname="Natalia" lastname="Chestkowska" birthdate="2006-10-01" gender="F" nation="POL" license="104115600047" swrid="5249565" athleteid="1895">
              <RESULTS>
                <RESULT eventid="1071" points="285" reactiontime="+84" swimtime="00:00:35.93" resultid="1896" heatid="2954" lane="6" entrytime="00:00:35.91" entrycourse="LCM" />
                <RESULT eventid="1111" points="296" reactiontime="+75" swimtime="00:01:36.19" resultid="1897" heatid="3004" lane="0" entrytime="00:01:35.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="265" reactiontime="+78" swimtime="00:01:20.46" resultid="1898" heatid="3030" lane="6" entrytime="00:01:21.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="281" reactiontime="+83" swimtime="00:00:44.87" resultid="1899" heatid="3047" lane="4" entrytime="00:00:43.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Janiak" birthdate="2008-03-01" gender="F" nation="POL" license="104115600087" swrid="5214625" athleteid="1921">
              <RESULTS>
                <RESULT eventid="1071" points="343" reactiontime="+66" swimtime="00:00:33.79" resultid="1922" heatid="2954" lane="9" />
                <RESULT eventid="1095" points="322" swimtime="00:00:39.36" resultid="1923" heatid="2984" lane="5" />
                <RESULT eventid="1119" points="307" swimtime="00:00:36.18" resultid="1924" heatid="3013" lane="2" />
                <RESULT eventid="1135" points="300" swimtime="00:01:17.18" resultid="1925" heatid="3029" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="214" swimtime="00:00:49.09" resultid="1926" heatid="3046" lane="5" />
                <RESULT eventid="1167" points="279" swimtime="00:03:12.95" resultid="1927" heatid="3066" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                    <SPLIT distance="100" swimtime="00:01:30.42" />
                    <SPLIT distance="150" swimtime="00:02:32.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kornelia" lastname="Salzman" birthdate="2010-07-23" gender="F" nation="POL" license="104115600178" swrid="5448040" athleteid="1944">
              <RESULTS>
                <RESULT eventid="1087" points="137" reactiontime="+61" swimtime="00:01:47.60" resultid="1945" heatid="2977" lane="5" entrytime="00:01:47.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="188" reactiontime="+75" swimtime="00:00:42.59" resultid="1946" heatid="3014" lane="9" entrytime="00:00:42.64" entrycourse="LCM" />
                <RESULT eventid="1135" points="215" reactiontime="+69" swimtime="00:01:26.26" resultid="1947" heatid="3029" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Klaudia" lastname="Borkiewicz" birthdate="2006-07-21" gender="F" nation="POL" license="104115600034" swrid="5009625" athleteid="1889">
              <RESULTS>
                <RESULT eventid="1071" points="547" reactiontime="+77" swimtime="00:00:28.94" resultid="1890" heatid="2959" lane="9" entrytime="00:00:28.38" entrycourse="LCM" />
                <RESULT comment="G2 - Pływak zanurzył się całkowicie w trakcie wyścigu (z wyjątkiem 15 m po starcie lub nawrocie)." eventid="1095" reactiontime="+67" status="DSQ" swimtime="00:00:00.00" resultid="1891" heatid="2987" lane="6" entrytime="00:00:31.94" entrycourse="LCM" />
                <RESULT eventid="1119" points="518" reactiontime="+78" swimtime="00:00:30.40" resultid="1892" heatid="3016" lane="8" entrytime="00:00:30.04" entrycourse="LCM" />
                <RESULT eventid="1135" points="524" reactiontime="+72" swimtime="00:01:04.13" resultid="1893" heatid="3033" lane="8" entrytime="00:01:04.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="471" reactiontime="+71" swimtime="00:01:13.97" resultid="1894" heatid="3061" lane="4" entrytime="00:01:12.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Bidziński" birthdate="2006-06-28" gender="M" nation="POL" license="104115700040" swrid="5190174" athleteid="1928">
              <RESULTS>
                <RESULT eventid="1075" points="498" reactiontime="+72" swimtime="00:00:26.38" resultid="1929" heatid="2970" lane="7" entrytime="00:00:26.14" entrycourse="LCM" />
                <RESULT eventid="1099" points="413" reactiontime="+84" swimtime="00:00:32.21" resultid="1930" heatid="2992" lane="1" entrytime="00:00:31.91" entrycourse="LCM" />
                <RESULT eventid="1123" points="419" reactiontime="+81" swimtime="00:00:29.74" resultid="1931" heatid="3020" lane="6" />
                <RESULT eventid="1139" points="518" reactiontime="+48" swimtime="00:00:58.40" resultid="1932" heatid="3041" lane="5" entrytime="00:00:57.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Janiak" birthdate="2006-02-26" gender="F" nation="POL" license="104115600068" swrid="5197714" athleteid="1900">
              <RESULTS>
                <RESULT eventid="1071" points="479" reactiontime="+63" swimtime="00:00:30.24" resultid="1901" heatid="2957" lane="8" entrytime="00:00:30.05" entrycourse="LCM" />
                <RESULT eventid="1111" points="407" reactiontime="+55" swimtime="00:01:26.50" resultid="1902" heatid="3004" lane="5" entrytime="00:01:26.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="360" swimtime="00:00:34.34" resultid="1903" heatid="3014" lane="2" entrytime="00:00:34.53" entrycourse="LCM" />
                <RESULT eventid="1135" points="462" reactiontime="+68" swimtime="00:01:06.87" resultid="1904" heatid="3032" lane="6" entrytime="00:01:07.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="417" reactiontime="+67" swimtime="00:00:39.35" resultid="1905" heatid="3048" lane="7" entrytime="00:00:39.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwier" lastname="Andrzejewski" birthdate="2009-02-09" gender="M" nation="POL" license="104115700160" swrid="5322504" athleteid="1933">
              <RESULTS>
                <RESULT eventid="1075" points="249" reactiontime="+80" swimtime="00:00:33.23" resultid="1934" heatid="2962" lane="2" />
                <RESULT eventid="1115" points="165" swimtime="00:01:43.69" resultid="1935" heatid="3007" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="129" reactiontime="+70" swimtime="00:00:43.97" resultid="1936" heatid="3018" lane="6" />
                <RESULT eventid="1139" points="250" reactiontime="+65" swimtime="00:01:14.43" resultid="1937" heatid="3037" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="201" reactiontime="+68" swimtime="00:00:44.30" resultid="1938" heatid="3050" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Grabiński" birthdate="2009-01-02" gender="M" nation="POL" license="104115700176" swrid="5322582" athleteid="1939">
              <RESULTS>
                <RESULT eventid="1075" points="206" reactiontime="+91" swimtime="00:00:35.37" resultid="1940" heatid="2963" lane="5" />
                <RESULT eventid="1115" points="207" reactiontime="+74" swimtime="00:01:36.13" resultid="1941" heatid="3006" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="201" reactiontime="+86" swimtime="00:01:20.01" resultid="1942" heatid="3036" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="213" reactiontime="+69" swimtime="00:00:43.40" resultid="1943" heatid="3052" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Zielińska" birthdate="2009-01-18" gender="F" nation="POL" license="104115600145" swrid="5322539" athleteid="1911">
              <RESULTS>
                <RESULT eventid="1071" points="348" swimtime="00:00:33.64" resultid="1912" heatid="2953" lane="2" />
                <RESULT eventid="1095" points="255" reactiontime="+95" swimtime="00:00:42.54" resultid="1913" heatid="2985" lane="7" />
                <RESULT eventid="1111" points="260" reactiontime="+84" swimtime="00:01:40.43" resultid="1914" heatid="3003" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="324" reactiontime="+82" swimtime="00:00:42.79" resultid="1915" heatid="3044" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Janiak" birthdate="2010-01-18" gender="F" nation="POL" license="104115600126" swrid="5271535" athleteid="1906">
              <RESULTS>
                <RESULT eventid="1071" points="287" swimtime="00:00:35.87" resultid="1907" heatid="2951" lane="7" />
                <RESULT eventid="1095" points="251" reactiontime="+56" swimtime="00:00:42.77" resultid="1908" heatid="2983" lane="5" />
                <RESULT eventid="1119" points="153" swimtime="00:00:45.59" resultid="1909" heatid="3012" lane="7" />
                <RESULT eventid="1159" points="227" reactiontime="+63" swimtime="00:01:34.32" resultid="1910" heatid="3060" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Chestkowska" birthdate="2009-05-12" gender="F" nation="POL" license="104115600048" swrid="5249566" athleteid="1948">
              <RESULTS>
                <RESULT eventid="1095" points="341" reactiontime="+70" swimtime="00:00:38.60" resultid="1949" heatid="2985" lane="1" />
                <RESULT eventid="1119" points="234" swimtime="00:00:39.60" resultid="1950" heatid="3013" lane="9" />
                <RESULT eventid="1143" points="299" reactiontime="+69" swimtime="00:00:43.94" resultid="1951" heatid="3045" lane="3" />
                <RESULT eventid="1159" points="297" reactiontime="+74" swimtime="00:01:26.22" resultid="1952" heatid="3060" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Krawczyk" birthdate="2008-09-23" gender="F" nation="POL" license="104115600117" swrid="5311268" athleteid="1953">
              <RESULTS>
                <RESULT eventid="1095" points="264" reactiontime="+75" swimtime="00:00:42.04" resultid="1954" heatid="2985" lane="4" entrytime="00:00:43.18" entrycourse="LCM" />
                <RESULT eventid="1119" points="181" reactiontime="+70" swimtime="00:00:43.17" resultid="1955" heatid="3014" lane="0" entrytime="00:00:41.72" entrycourse="LCM" />
                <RESULT eventid="1135" points="225" reactiontime="+72" swimtime="00:01:24.98" resultid="1956" heatid="3029" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="211" reactiontime="+76" swimtime="00:03:31.54" resultid="1957" heatid="3067" lane="3" entrytime="00:03:31.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                    <SPLIT distance="100" swimtime="00:01:38.58" />
                    <SPLIT distance="150" swimtime="00:02:42.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Cicha" birthdate="2008-11-07" gender="F" nation="POL" license="104115600109" swrid="5322568" athleteid="1916">
              <RESULTS>
                <RESULT eventid="1071" points="311" reactiontime="+82" swimtime="00:00:34.90" resultid="1917" heatid="2951" lane="3" />
                <RESULT eventid="1095" points="353" reactiontime="+82" swimtime="00:00:38.15" resultid="1918" heatid="2985" lane="8" />
                <RESULT eventid="1119" points="251" reactiontime="+77" swimtime="00:00:38.71" resultid="1919" heatid="3012" lane="2" />
                <RESULT eventid="1143" points="212" swimtime="00:00:49.30" resultid="1920" heatid="3046" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+77" swimtime="00:02:00.08" resultid="1958" heatid="2948" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="100" swimtime="00:01:04.77" />
                    <SPLIT distance="150" swimtime="00:01:34.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1889" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="1895" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="1900" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="1928" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1183" reactiontime="+64" swimtime="00:02:17.27" resultid="1959" heatid="3079" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="150" swimtime="00:01:50.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1889" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="1895" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="1900" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="1928" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1183" reactiontime="+77" swimtime="00:02:36.63" resultid="1960" heatid="3079" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                    <SPLIT distance="100" swimtime="00:01:22.38" />
                    <SPLIT distance="150" swimtime="00:02:01.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1948" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="1911" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="1916" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="1921" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="07911" nation="POL" region="11" clubid="2419" name="Uks &quot;Via Sport&quot;">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Kapka" birthdate="1977-11-05" gender="M" nation="POL" license="107911700092" athleteid="2420">
              <RESULTS>
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie)." eventid="1083" reactiontime="+87" status="DSQ" swimtime="00:00:00.00" resultid="2421" heatid="2975" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:01:33.73" />
                    <SPLIT distance="150" swimtime="00:02:27.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="233" reactiontime="+76" swimtime="00:01:32.36" resultid="2422" heatid="3007" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="189" reactiontime="+79" swimtime="00:03:14.88" resultid="2423" heatid="3027" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.02" />
                    <SPLIT distance="100" swimtime="00:01:37.32" />
                    <SPLIT distance="150" swimtime="00:02:28.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="2424" heatid="3063" lane="5" />
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="2425" heatid="3070" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00402" nation="POL" region="02" clubid="2449" name="UKS ,,Ósemka&apos;&apos; Toruń">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Jackiewicz" birthdate="2008-02-21" gender="F" nation="POL" license="100402600058" swrid="5108151" athleteid="2450">
              <RESULTS>
                <RESULT eventid="1071" points="470" reactiontime="+62" swimtime="00:00:30.43" resultid="2451" heatid="2956" lane="5" entrytime="00:00:30.20" entrycourse="LCM" />
                <RESULT eventid="1087" points="350" reactiontime="+70" swimtime="00:01:18.69" resultid="2452" heatid="2978" lane="0" entrytime="00:01:18.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="387" reactiontime="+70" swimtime="00:00:33.50" resultid="2453" heatid="3015" lane="0" entrytime="00:00:32.67" entrycourse="LCM" />
                <RESULT eventid="1143" points="378" reactiontime="+63" swimtime="00:00:40.63" resultid="2454" heatid="3046" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="501713" nation="POL" region="13" clubid="2809" name="TP Masters Olsztyn">
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Sokulski" birthdate="1991-02-10" gender="M" nation="POL" license="101713700005" swrid="4062177" athleteid="2805">
              <RESULTS>
                <RESULT eventid="1075" points="645" reactiontime="+69" swimtime="00:00:24.19" resultid="2806" heatid="2971" lane="5" entrytime="00:00:23.99" entrycourse="LCM" />
                <RESULT eventid="1123" points="666" reactiontime="+70" swimtime="00:00:25.49" resultid="2807" heatid="3024" lane="3" entrytime="00:00:25.06" entrycourse="LCM" />
                <RESULT eventid="1139" points="662" reactiontime="+67" swimtime="00:00:53.81" resultid="2808" heatid="3036" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01014" nation="POL" region="14" clubid="1362" name="KS ,,1&apos;&apos; Ożarów Mazowiecki">
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Popow" birthdate="2006-04-09" gender="M" nation="POL" license="101014700117" swrid="5161556" athleteid="1374">
              <RESULTS>
                <RESULT eventid="1099" status="DNS" swimtime="00:00:00.00" resultid="1375" heatid="2993" lane="7" entrytime="00:00:29.11" entrycourse="LCM" />
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="1376" heatid="3001" lane="8" entrytime="00:02:09.59" entrycourse="LCM" />
                <RESULT eventid="1131" status="DNS" swimtime="00:00:00.00" resultid="1377" heatid="3028" lane="5" entrytime="00:02:17.59" entrycourse="LCM" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="1378" heatid="3065" lane="5" entrytime="00:01:02.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Gajda" birthdate="2006-09-08" gender="F" nation="POL" license="101014600116" swrid="5161565" athleteid="1363">
              <RESULTS>
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="1364" heatid="2958" lane="1" entrytime="00:00:28.86" entrycourse="LCM" />
                <RESULT eventid="1095" status="DNS" swimtime="00:00:00.00" resultid="1365" heatid="2986" lane="6" entrytime="00:00:35.53" entrycourse="LCM" />
                <RESULT eventid="1135" status="DNS" swimtime="00:00:00.00" resultid="1366" heatid="3033" lane="7" entrytime="00:01:04.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Adamczyk" birthdate="2006-04-28" gender="F" nation="POL" license="101014600111" swrid="5056861" athleteid="1369">
              <RESULTS>
                <RESULT eventid="1087" status="DNS" swimtime="00:00:00.00" resultid="1370" heatid="2979" lane="8" entrytime="00:01:08.07" entrycourse="LCM" />
                <RESULT eventid="1103" status="DNS" swimtime="00:00:00.00" resultid="1371" heatid="2997" lane="2" entrytime="00:02:14.60" entrycourse="LCM" />
                <RESULT eventid="1119" status="DNS" swimtime="00:00:00.00" resultid="1372" heatid="3015" lane="6" entrytime="00:00:31.19" entrycourse="LCM" />
                <RESULT eventid="1135" status="DNS" swimtime="00:00:00.00" resultid="1373" heatid="3034" lane="9" entrytime="00:01:02.13" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Liszkiewicz" birthdate="2006-04-30" gender="M" nation="POL" license="101014700127" swrid="5331237" athleteid="1367">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="1368" heatid="2960" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="1379" heatid="2948" lane="0" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02302" nation="POL" region="02" clubid="2444" name="Uks ,,Orka&apos;&apos; Mogilno">
          <ATHLETES>
            <ATHLETE firstname="Weronika" lastname="Michalska" birthdate="2006-03-31" gender="F" nation="POL" license="102302600005" swrid="5114182" athleteid="2445">
              <RESULTS>
                <RESULT eventid="1071" points="525" reactiontime="+80" swimtime="00:00:29.33" resultid="2446" heatid="2957" lane="3" entrytime="00:00:29.48" entrycourse="LCM" />
                <RESULT eventid="1095" points="541" reactiontime="+66" swimtime="00:00:33.11" resultid="2447" heatid="2987" lane="8" entrytime="00:00:32.42" entrycourse="LCM" />
                <RESULT eventid="1119" points="461" reactiontime="+74" swimtime="00:00:31.62" resultid="2448" heatid="3015" lane="1" entrytime="00:00:31.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01015" nation="POL" region="15" clubid="2686" name="UKS Trójka Środa Wlkp.">
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Kucharska" birthdate="2005-01-04" gender="F" nation="POL" license="101015600037" swrid="5096958" athleteid="2697">
              <RESULTS>
                <RESULT eventid="1071" points="571" swimtime="00:00:28.53" resultid="2698" heatid="2951" lane="2" />
                <RESULT eventid="1111" points="481" reactiontime="+68" swimtime="00:01:21.82" resultid="2699" heatid="3005" lane="1" entrytime="00:01:19.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="542" reactiontime="+77" swimtime="00:01:03.42" resultid="2700" heatid="3030" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="609" reactiontime="+65" swimtime="00:00:34.68" resultid="2701" heatid="3049" lane="5" entrytime="00:00:34.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Waleron" birthdate="2010-04-06" gender="M" nation="POL" license="101015700078" swrid="5448042" athleteid="2712">
              <RESULTS>
                <RESULT eventid="1091" points="118" swimtime="00:01:40.70" resultid="2713" heatid="2980" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="142" reactiontime="+65" swimtime="00:01:48.84" resultid="2714" heatid="3006" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="120" reactiontime="+67" swimtime="00:00:45.07" resultid="2715" heatid="3018" lane="1" />
                <RESULT eventid="1147" points="138" swimtime="00:00:50.14" resultid="2716" heatid="3051" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelina" lastname="Mieloch" birthdate="2005-07-24" gender="F" nation="POL" license="101015600044" swrid="5117134" athleteid="2702">
              <RESULTS>
                <RESULT eventid="1071" points="473" reactiontime="+63" swimtime="00:00:30.37" resultid="2703" heatid="2952" lane="4" />
                <RESULT eventid="1095" points="433" reactiontime="+65" swimtime="00:00:35.66" resultid="2704" heatid="2986" lane="5" entrytime="00:00:35.14" entrycourse="LCM" />
                <RESULT eventid="1127" points="375" reactiontime="+66" swimtime="00:02:51.00" resultid="2705" heatid="3026" lane="2" entrytime="00:02:50.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:22.48" />
                    <SPLIT distance="150" swimtime="00:02:07.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="378" reactiontime="+66" swimtime="00:01:19.62" resultid="2706" heatid="3061" lane="5" entrytime="00:01:16.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Nowak" birthdate="2005-08-04" gender="M" nation="POL" license="101015700036" swrid="5117131" athleteid="2707">
              <RESULTS>
                <RESULT eventid="1075" points="470" reactiontime="+82" swimtime="00:00:26.89" resultid="2708" heatid="2969" lane="8" entrytime="00:00:27.23" entrycourse="LCM" />
                <RESULT eventid="1091" points="403" reactiontime="+61" swimtime="00:01:06.99" resultid="2709" heatid="2981" lane="5" entrytime="00:01:07.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="449" reactiontime="+73" swimtime="00:00:29.08" resultid="2710" heatid="3022" lane="6" entrytime="00:00:29.51" entrycourse="LCM" />
                <RESULT eventid="1139" points="503" reactiontime="+73" swimtime="00:00:58.97" resultid="2711" heatid="3041" lane="8" entrytime="00:00:59.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Perlik" birthdate="2006-09-24" gender="F" nation="POL" license="101015600057" swrid="5153534" athleteid="2692">
              <RESULTS>
                <RESULT eventid="1071" points="480" reactiontime="+85" swimtime="00:00:30.23" resultid="2693" heatid="2957" lane="9" entrytime="00:00:30.05" entrycourse="LCM" />
                <RESULT eventid="1087" points="372" reactiontime="+85" swimtime="00:01:17.09" resultid="2694" heatid="2978" lane="8" entrytime="00:01:17.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="406" reactiontime="+81" swimtime="00:00:32.97" resultid="2695" heatid="3014" lane="4" entrytime="00:00:33.80" entrycourse="LCM" />
                <RESULT eventid="1135" points="432" reactiontime="+80" swimtime="00:01:08.38" resultid="2696" heatid="3033" lane="9" entrytime="00:01:06.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Waleron" birthdate="2008-09-11" gender="M" nation="POL" license="101015700077" swrid="5334854" athleteid="2687">
              <RESULTS>
                <RESULT eventid="1067" points="228" swimtime="00:06:38.89" resultid="2688" heatid="2950" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                    <SPLIT distance="100" swimtime="00:01:35.81" />
                    <SPLIT distance="150" swimtime="00:02:25.89" />
                    <SPLIT distance="200" swimtime="00:03:14.78" />
                    <SPLIT distance="250" swimtime="00:04:12.18" />
                    <SPLIT distance="300" swimtime="00:05:09.03" />
                    <SPLIT distance="350" swimtime="00:05:55.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="222" reactiontime="+80" swimtime="00:00:39.59" resultid="2689" heatid="2990" lane="7" />
                <RESULT eventid="1107" points="230" swimtime="00:02:46.37" resultid="2690" heatid="2998" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                    <SPLIT distance="100" swimtime="00:01:22.30" />
                    <SPLIT distance="150" swimtime="00:02:05.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="217" reactiontime="+77" swimtime="00:03:06.04" resultid="2691" heatid="3027" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.75" />
                    <SPLIT distance="100" swimtime="00:01:33.18" />
                    <SPLIT distance="150" swimtime="00:02:21.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00802" nation="POL" region="02" clubid="2230" name="MUKS &apos;&apos;Piętnastka&apos;&apos;">
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Sobieralski" birthdate="2008-11-26" gender="M" nation="POL" license="100802700252" swrid="5350180" athleteid="2284">
              <RESULTS>
                <RESULT eventid="1075" points="341" reactiontime="+77" swimtime="00:00:29.92" resultid="2285" heatid="2967" lane="5" entrytime="00:00:29.54" entrycourse="LCM" />
                <RESULT eventid="1099" points="298" reactiontime="+74" swimtime="00:00:35.91" resultid="2286" heatid="2991" lane="3" entrytime="00:00:35.59" entrycourse="LCM" />
                <RESULT eventid="1123" points="308" reactiontime="+77" swimtime="00:00:32.97" resultid="2287" heatid="3021" lane="6" entrytime="00:00:32.73" entrycourse="LCM" />
                <RESULT eventid="1147" points="253" reactiontime="+75" swimtime="00:00:40.98" resultid="2288" heatid="3055" lane="6" entrytime="00:00:40.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Melissa" lastname="Orum" birthdate="2004-09-17" gender="F" nation="POL" license="100802600197" swrid="5075949" athleteid="2270">
              <RESULTS>
                <RESULT eventid="1071" points="531" swimtime="00:00:29.22" resultid="2271" heatid="2958" lane="2" entrytime="00:00:28.75" entrycourse="LCM" />
                <RESULT eventid="1103" points="511" reactiontime="+78" swimtime="00:02:21.28" resultid="2272" heatid="2994" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                    <SPLIT distance="150" swimtime="00:01:45.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="443" reactiontime="+75" swimtime="00:00:38.55" resultid="2273" heatid="3045" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Kowalczyk" birthdate="2008-03-24" gender="M" nation="POL" license="100802700203" swrid="5087091" athleteid="2245">
              <RESULTS>
                <RESULT eventid="1067" points="336" reactiontime="+67" swimtime="00:05:50.63" resultid="2246" heatid="2950" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:20.54" />
                    <SPLIT distance="150" swimtime="00:02:04.64" />
                    <SPLIT distance="200" swimtime="00:02:47.61" />
                    <SPLIT distance="250" swimtime="00:03:36.76" />
                    <SPLIT distance="300" swimtime="00:04:26.86" />
                    <SPLIT distance="350" swimtime="00:05:09.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="321" swimtime="00:03:04.12" resultid="2247" heatid="2974" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:01:30.90" />
                    <SPLIT distance="150" swimtime="00:02:18.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="311" swimtime="00:02:30.46" resultid="2248" heatid="3000" lane="1" entrytime="00:02:26.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:53.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="362" reactiontime="+69" swimtime="00:02:36.98" resultid="2249" heatid="3027" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                    <SPLIT distance="100" swimtime="00:01:17.54" />
                    <SPLIT distance="150" swimtime="00:01:58.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="338" reactiontime="+55" swimtime="00:02:43.60" resultid="2250" heatid="3072" lane="9" entrytime="00:02:40.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                    <SPLIT distance="100" swimtime="00:01:17.35" />
                    <SPLIT distance="150" swimtime="00:02:04.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Woroniecka" birthdate="2005-02-19" gender="F" nation="POL" license="100802600231" swrid="4907608" athleteid="2326">
              <RESULTS>
                <RESULT eventid="1095" points="494" reactiontime="+79" swimtime="00:00:34.12" resultid="2327" heatid="2983" lane="4" />
                <RESULT eventid="1103" points="514" reactiontime="+84" swimtime="00:02:20.96" resultid="2328" heatid="2996" lane="6" entrytime="00:02:25.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:07.60" />
                    <SPLIT distance="150" swimtime="00:01:43.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="533" reactiontime="+79" swimtime="00:01:03.75" resultid="2329" heatid="3033" lane="1" entrytime="00:01:04.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matylda" lastname="Antkowiak" birthdate="2007-01-17" gender="F" nation="POL" license="100802600312" swrid="5264076" athleteid="2266">
              <RESULTS>
                <RESULT eventid="1071" points="363" reactiontime="+92" swimtime="00:00:33.16" resultid="2267" heatid="2955" lane="7" entrytime="00:00:32.71" entrycourse="LCM" />
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="2268" heatid="3003" lane="3" />
                <RESULT eventid="1135" points="391" reactiontime="+53" swimtime="00:01:10.68" resultid="2269" heatid="3031" lane="5" entrytime="00:01:10.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Nowak" birthdate="2005-07-02" gender="F" nation="POL" license="100802600311" swrid="4943255" athleteid="2301">
              <RESULTS>
                <RESULT eventid="1087" points="489" reactiontime="+52" swimtime="00:01:10.38" resultid="2302" heatid="2978" lane="5" entrytime="00:01:08.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="486" reactiontime="+44" swimtime="00:00:31.07" resultid="2303" heatid="3015" lane="5" entrytime="00:00:30.60" entrycourse="LCM" />
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="2304" heatid="3074" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Ronkiewicz" birthdate="2005-01-17" gender="F" nation="POL" license="100802600218" swrid="4756930" athleteid="2351">
              <RESULTS>
                <RESULT eventid="1119" points="432" reactiontime="+75" swimtime="00:00:32.30" resultid="2352" heatid="3011" lane="3" />
                <RESULT eventid="1143" points="545" reactiontime="+68" swimtime="00:00:35.98" resultid="2353" heatid="3049" lane="2" entrytime="00:00:35.45" entrycourse="LCM" />
                <RESULT eventid="1167" points="488" reactiontime="+74" swimtime="00:02:40.12" resultid="2354" heatid="3066" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                    <SPLIT distance="100" swimtime="00:01:16.25" />
                    <SPLIT distance="150" swimtime="00:02:02.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Matjakowska" birthdate="2006-04-09" gender="F" nation="POL" license="100802600281" swrid="4990961" athleteid="2297">
              <RESULTS>
                <RESULT eventid="1087" points="339" reactiontime="+79" swimtime="00:01:19.53" resultid="2298" heatid="2977" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="404" reactiontime="+80" swimtime="00:00:36.48" resultid="2299" heatid="2984" lane="3" />
                <RESULT eventid="1119" points="354" reactiontime="+75" swimtime="00:00:34.52" resultid="2300" heatid="3012" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pola" lastname="Karolczak" birthdate="2006-04-13" gender="F" nation="POL" license="100802600286" swrid="5112761" athleteid="2241">
              <RESULTS>
                <RESULT eventid="1063" points="464" reactiontime="+83" swimtime="00:05:43.89" resultid="2242" heatid="2949" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:16.55" />
                    <SPLIT distance="150" swimtime="00:02:00.88" />
                    <SPLIT distance="200" swimtime="00:02:44.56" />
                    <SPLIT distance="250" swimtime="00:03:32.02" />
                    <SPLIT distance="300" swimtime="00:04:21.44" />
                    <SPLIT distance="350" swimtime="00:05:02.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="484" reactiontime="+76" swimtime="00:00:34.34" resultid="2243" heatid="2984" lane="2" />
                <RESULT eventid="1119" points="458" reactiontime="+77" swimtime="00:00:31.68" resultid="2244" heatid="3013" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojtek" lastname="Sobieralski" birthdate="2010-12-21" gender="M" nation="POL" license="100802700355" swrid="5460449" athleteid="2279">
              <RESULTS>
                <RESULT eventid="1075" points="162" reactiontime="+101" swimtime="00:00:38.28" resultid="2280" heatid="2965" lane="2" entrytime="00:00:39.60" entrycourse="LCM" />
                <RESULT eventid="1099" points="108" reactiontime="+99" swimtime="00:00:50.31" resultid="2281" heatid="2990" lane="4" entrytime="00:00:47.78" entrycourse="LCM" />
                <RESULT eventid="1123" points="68" reactiontime="+94" swimtime="00:00:54.55" resultid="2282" heatid="3021" lane="0" entrytime="00:00:49.47" entrycourse="LCM" />
                <RESULT eventid="1163" points="102" reactiontime="+79" swimtime="00:01:50.88" resultid="2283" heatid="3064" lane="8" entrytime="00:01:46.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Jaworska" birthdate="2005-07-22" gender="F" nation="POL" license="100802600243" swrid="5056997" athleteid="2274">
              <RESULTS>
                <RESULT eventid="1071" points="467" reactiontime="+78" swimtime="00:00:30.49" resultid="2275" heatid="2952" lane="5" />
                <RESULT eventid="1119" points="422" reactiontime="+75" swimtime="00:00:32.57" resultid="2276" heatid="3013" lane="7" />
                <RESULT eventid="1135" points="502" reactiontime="+77" swimtime="00:01:05.05" resultid="2277" heatid="3032" lane="4" entrytime="00:01:06.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="466" reactiontime="+59" swimtime="00:02:42.57" resultid="2278" heatid="3066" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:16.42" />
                    <SPLIT distance="150" swimtime="00:02:06.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adriana" lastname="Kulczyńska" birthdate="2006-10-12" gender="F" nation="POL" license="100802600237" swrid="4907680" athleteid="2322">
              <RESULTS>
                <RESULT eventid="1095" points="483" reactiontime="+69" swimtime="00:00:34.38" resultid="2323" heatid="2986" lane="2" entrytime="00:00:35.60" entrycourse="LCM" />
                <RESULT eventid="1127" points="470" reactiontime="+66" swimtime="00:02:38.55" resultid="2324" heatid="3026" lane="3" entrytime="00:02:39.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:14.36" />
                    <SPLIT distance="150" swimtime="00:01:57.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="465" reactiontime="+78" swimtime="00:02:42.73" resultid="2325" heatid="3068" lane="7" entrytime="00:02:47.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="150" swimtime="00:02:03.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Knopp" birthdate="2004-06-22" gender="M" nation="POL" license="100802700200" swrid="4907694" athleteid="2309">
              <RESULTS>
                <RESULT eventid="1091" points="552" reactiontime="+73" swimtime="00:01:00.33" resultid="2310" heatid="2982" lane="6" entrytime="00:00:59.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="511" reactiontime="+84" swimtime="00:00:27.85" resultid="2311" heatid="3020" lane="9" />
                <RESULT eventid="1155" points="528" reactiontime="+72" swimtime="00:02:16.93" resultid="2312" heatid="3059" lane="4" entrytime="00:02:15.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                    <SPLIT distance="100" swimtime="00:01:05.97" />
                    <SPLIT distance="150" swimtime="00:01:42.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelina" lastname="Moritz" birthdate="2005-09-15" gender="F" nation="POL" license="100802600229" swrid="4907603" athleteid="2337">
              <RESULTS>
                <RESULT eventid="1103" points="522" reactiontime="+83" swimtime="00:02:20.28" resultid="2338" heatid="2997" lane="9" entrytime="00:02:20.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:06.54" />
                    <SPLIT distance="150" swimtime="00:01:43.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="371" reactiontime="+82" swimtime="00:00:33.98" resultid="2339" heatid="3012" lane="9" />
                <RESULT eventid="1135" points="489" reactiontime="+73" swimtime="00:01:05.62" resultid="2340" heatid="3029" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="454" swimtime="00:02:44.05" resultid="2341" heatid="3068" lane="2" entrytime="00:02:37.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:02:05.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Janeczek" birthdate="2004-06-01" gender="M" nation="POL" license="100802700212" swrid="4907622" athleteid="2294">
              <RESULTS>
                <RESULT eventid="1083" points="494" reactiontime="+79" swimtime="00:02:39.47" resultid="2295" heatid="2975" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                    <SPLIT distance="150" swimtime="00:01:57.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="513" swimtime="00:02:22.32" resultid="2296" heatid="3070" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                    <SPLIT distance="100" swimtime="00:01:07.06" />
                    <SPLIT distance="150" swimtime="00:01:48.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Sędłak" birthdate="2005-01-17" gender="F" nation="POL" license="100802600221" swrid="4980030" athleteid="2236">
              <RESULTS>
                <RESULT eventid="1063" points="590" reactiontime="+76" swimtime="00:05:17.54" resultid="2237" heatid="2949" lane="4" entrytime="00:05:20.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:10.29" />
                    <SPLIT distance="150" swimtime="00:01:50.76" />
                    <SPLIT distance="200" swimtime="00:02:31.78" />
                    <SPLIT distance="250" swimtime="00:03:15.62" />
                    <SPLIT distance="300" swimtime="00:04:01.91" />
                    <SPLIT distance="350" swimtime="00:04:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="563" reactiontime="+69" swimtime="00:00:29.57" resultid="2238" heatid="3012" lane="6" />
                <RESULT eventid="1143" points="582" reactiontime="+69" swimtime="00:00:35.20" resultid="2239" heatid="3044" lane="3" />
                <RESULT eventid="1167" points="615" reactiontime="+74" swimtime="00:02:28.23" resultid="2240" heatid="3068" lane="4" entrytime="00:02:27.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:11.49" />
                    <SPLIT distance="150" swimtime="00:01:53.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Pasik" birthdate="2007-01-28" gender="F" nation="POL" license="100802600292" swrid="4997805" athleteid="2313">
              <RESULTS>
                <RESULT eventid="1095" points="311" reactiontime="+72" swimtime="00:00:39.80" resultid="2314" heatid="2985" lane="6" />
                <RESULT eventid="1103" points="294" reactiontime="+78" swimtime="00:02:49.73" resultid="2315" heatid="2995" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:19.76" />
                    <SPLIT distance="150" swimtime="00:02:04.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="325" reactiontime="+69" swimtime="00:02:59.31" resultid="2316" heatid="3025" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                    <SPLIT distance="100" swimtime="00:01:26.18" />
                    <SPLIT distance="150" swimtime="00:02:12.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="341" reactiontime="+67" swimtime="00:00:42.08" resultid="2317" heatid="3046" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Miniszewski" birthdate="2004-01-31" gender="M" nation="POL" license="100802700199" swrid="5027959" athleteid="2342">
              <RESULTS>
                <RESULT eventid="1107" points="574" reactiontime="+66" swimtime="00:02:02.72" resultid="2343" heatid="3001" lane="5" entrytime="00:02:02.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                    <SPLIT distance="100" swimtime="00:01:00.03" />
                    <SPLIT distance="150" swimtime="00:01:31.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="620" reactiontime="+70" swimtime="00:00:55.01" resultid="2344" heatid="3043" lane="6" entrytime="00:00:54.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="489" reactiontime="+69" swimtime="00:02:20.47" resultid="2345" heatid="3059" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                    <SPLIT distance="100" swimtime="00:01:05.05" />
                    <SPLIT distance="150" swimtime="00:01:41.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Brucka" birthdate="2006-07-11" gender="F" nation="POL" license="100802600279" swrid="4990960" athleteid="2330">
              <RESULTS>
                <RESULT eventid="1095" points="385" reactiontime="+70" swimtime="00:00:37.06" resultid="2331" heatid="2984" lane="8" />
                <RESULT eventid="1119" points="380" reactiontime="+64" swimtime="00:00:33.71" resultid="2332" heatid="3012" lane="8" />
                <RESULT eventid="1167" points="407" reactiontime="+63" swimtime="00:02:50.05" resultid="2333" heatid="3067" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:20.55" />
                    <SPLIT distance="150" swimtime="00:02:11.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Rostkowski" birthdate="2006-04-22" gender="M" nation="POL" license="100802700284" swrid="5056999" athleteid="2305">
              <RESULTS>
                <RESULT eventid="1091" points="407" reactiontime="+79" swimtime="00:01:06.77" resultid="2306" heatid="2982" lane="9" entrytime="00:01:05.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="431" reactiontime="+73" swimtime="00:00:29.47" resultid="2307" heatid="3018" lane="2" />
                <RESULT eventid="1163" points="369" reactiontime="+67" swimtime="00:01:12.26" resultid="2308" heatid="3064" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Hermanowska" birthdate="2004-12-15" gender="F" nation="POL" license="100802600202" swrid="4907692" athleteid="2318">
              <RESULTS>
                <RESULT eventid="1095" points="543" reactiontime="+76" swimtime="00:00:33.06" resultid="2319" heatid="2985" lane="2" />
                <RESULT eventid="1111" points="562" reactiontime="+75" swimtime="00:01:17.67" resultid="2320" heatid="3005" lane="5" entrytime="00:01:14.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="617" reactiontime="+72" swimtime="00:00:34.52" resultid="2321" heatid="3049" lane="4" entrytime="00:00:33.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Pytloch" birthdate="2005-10-29" gender="F" nation="POL" license="100802600309" swrid="4928417" athleteid="2260">
              <RESULTS>
                <RESULT eventid="1071" points="564" reactiontime="+69" swimtime="00:00:28.64" resultid="2261" heatid="2958" lane="0" entrytime="00:00:28.91" entrycourse="LCM" />
                <RESULT eventid="1087" points="542" swimtime="00:01:08.04" resultid="2262" heatid="2979" lane="2" entrytime="00:01:06.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="508" reactiontime="+70" swimtime="00:00:30.61" resultid="2263" heatid="3015" lane="4" entrytime="00:00:30.32" entrycourse="LCM" />
                <RESULT eventid="1135" points="566" reactiontime="+67" swimtime="00:01:02.48" resultid="2264" heatid="3030" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="524" reactiontime="+67" swimtime="00:02:36.40" resultid="2265" heatid="3067" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:16.29" />
                    <SPLIT distance="150" swimtime="00:02:02.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Bania" birthdate="2005-09-10" gender="M" nation="POL" license="100802700219" swrid="5108576" athleteid="2251">
              <RESULTS>
                <RESULT eventid="1067" points="486" reactiontime="+76" swimtime="00:05:09.98" resultid="2252" heatid="2950" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:45.42" />
                    <SPLIT distance="200" swimtime="00:02:25.48" />
                    <SPLIT distance="250" swimtime="00:03:13.54" />
                    <SPLIT distance="300" swimtime="00:04:01.49" />
                    <SPLIT distance="350" swimtime="00:04:36.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="532" reactiontime="+81" swimtime="00:00:29.61" resultid="2253" heatid="2988" lane="3" />
                <RESULT eventid="1155" points="502" reactiontime="+70" swimtime="00:02:19.25" resultid="2254" heatid="3059" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="100" swimtime="00:01:06.28" />
                    <SPLIT distance="150" swimtime="00:01:43.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nadia" lastname="Studzińska" birthdate="2004-04-18" gender="F" nation="POL" license="100802600195" swrid="4001613" athleteid="2334">
              <RESULTS>
                <RESULT eventid="1103" points="484" reactiontime="+78" swimtime="00:02:23.86" resultid="2335" heatid="2995" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:08.76" />
                    <SPLIT distance="150" swimtime="00:01:46.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="452" reactiontime="+74" swimtime="00:01:14.99" resultid="2336" heatid="3061" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Sadowska" birthdate="2004-12-11" gender="F" nation="POL" license="100802600268" swrid="4907627" athleteid="2231">
              <RESULTS>
                <RESULT eventid="1063" points="492" reactiontime="+77" swimtime="00:05:37.39" resultid="2232" heatid="2949" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:11.74" />
                    <SPLIT distance="150" swimtime="00:01:55.57" />
                    <SPLIT distance="200" swimtime="00:02:37.89" />
                    <SPLIT distance="250" swimtime="00:03:27.48" />
                    <SPLIT distance="300" swimtime="00:04:19.41" />
                    <SPLIT distance="350" swimtime="00:04:58.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="458" reactiontime="+71" swimtime="00:00:34.98" resultid="2233" heatid="2985" lane="0" />
                <RESULT eventid="1135" points="559" reactiontime="+69" swimtime="00:01:02.76" resultid="2234" heatid="3033" lane="4" entrytime="00:01:02.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="467" reactiontime="+75" swimtime="00:02:36.91" resultid="2235" heatid="3058" lane="5" entrytime="00:02:39.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:14.02" />
                    <SPLIT distance="150" swimtime="00:01:55.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Szymański" birthdate="2005-01-09" gender="M" nation="POL" license="100802700220" swrid="4934162" athleteid="2255">
              <RESULTS>
                <RESULT eventid="1067" points="436" reactiontime="+75" swimtime="00:05:21.33" resultid="2256" heatid="2950" lane="5" entrytime="00:05:01.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:13.28" />
                    <SPLIT distance="150" swimtime="00:01:56.70" />
                    <SPLIT distance="200" swimtime="00:02:40.98" />
                    <SPLIT distance="250" swimtime="00:03:21.44" />
                    <SPLIT distance="300" swimtime="00:04:04.83" />
                    <SPLIT distance="350" swimtime="00:04:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie)." eventid="1083" reactiontime="+74" status="DSQ" swimtime="00:00:00.00" resultid="2257" heatid="2976" lane="3" entrytime="00:02:31.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="100" swimtime="00:01:13.12" />
                    <SPLIT distance="150" swimtime="00:01:53.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="545" reactiontime="+71" swimtime="00:01:09.63" resultid="2258" heatid="3010" lane="1" entrytime="00:01:09.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="531" reactiontime="+71" swimtime="00:02:20.76" resultid="2259" heatid="3070" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:09.65" />
                    <SPLIT distance="150" swimtime="00:01:48.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivier" lastname="Piątek" birthdate="2004-08-09" gender="M" nation="POL" license="100802700271" swrid="5027954" athleteid="2289">
              <RESULTS>
                <RESULT eventid="1075" points="578" reactiontime="+68" swimtime="00:00:25.10" resultid="2290" heatid="2971" lane="8" entrytime="00:00:24.99" entrycourse="LCM" />
                <RESULT eventid="1099" points="482" reactiontime="+68" swimtime="00:00:30.59" resultid="2291" heatid="2990" lane="0" />
                <RESULT eventid="1123" points="528" reactiontime="+70" swimtime="00:00:27.54" resultid="2292" heatid="3023" lane="3" entrytime="00:00:27.47" entrycourse="LCM" />
                <RESULT eventid="1147" points="480" reactiontime="+71" swimtime="00:00:33.14" resultid="2293" heatid="3052" lane="9" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+76" swimtime="00:01:57.14" resultid="2355" heatid="2948" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                    <SPLIT distance="100" swimtime="00:00:58.28" />
                    <SPLIT distance="150" swimtime="00:01:27.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2305" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="2245" number="2" reactiontime="+13" />
                    <RELAYPOSITION athleteid="2326" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="2337" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="O9 - Pływak niewłaściwie zachowywał się podczas zawodów (np. opóźnianie startu, umyślne zakłócanie porządku i inne)." eventid="1183" reactiontime="+63" status="DSQ" swimtime="00:00:00.00" resultid="2359" heatid="3079" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:06.50" />
                    <SPLIT distance="150" swimtime="00:01:33.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2270" number="1" reactiontime="+63" status="DSQ" />
                    <RELAYPOSITION athleteid="2318" number="2" reactiontime="+10" status="DSQ" />
                    <RELAYPOSITION athleteid="2289" number="3" reactiontime="+20" status="DSQ" />
                    <RELAYPOSITION athleteid="2294" number="4" reactiontime="+33" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+68" swimtime="00:01:45.45" resultid="2356" heatid="2948" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.92" />
                    <SPLIT distance="100" swimtime="00:00:49.60" />
                    <SPLIT distance="150" swimtime="00:01:16.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2289" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2294" number="2" />
                    <RELAYPOSITION athleteid="2318" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2270" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1183" reactiontime="+71" swimtime="00:02:00.17" resultid="2360" heatid="3079" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="100" swimtime="00:01:01.78" />
                    <SPLIT distance="150" swimtime="00:01:31.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2251" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="2255" number="2" />
                    <RELAYPOSITION athleteid="2236" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2260" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+80" swimtime="00:01:48.47" resultid="2357" heatid="2947" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.10" />
                    <SPLIT distance="100" swimtime="00:00:51.08" />
                    <SPLIT distance="150" swimtime="00:01:19.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2342" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2309" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="2231" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="2334" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1183" reactiontime="+71" swimtime="00:02:01.11" resultid="2361" heatid="3079" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:06.20" />
                    <SPLIT distance="150" swimtime="00:01:36.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2342" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="2334" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="2231" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2309" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+71" swimtime="00:01:50.01" resultid="2358" heatid="2948" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.29" />
                    <SPLIT distance="100" swimtime="00:00:52.70" />
                    <SPLIT distance="150" swimtime="00:01:21.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2251" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="2255" number="2" reactiontime="+24" />
                    <RELAYPOSITION athleteid="2301" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="2260" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1183" reactiontime="+66" swimtime="00:02:07.87" resultid="2362" heatid="3078" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:38.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2245" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2351" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="2305" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="2274" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="05415" nation="POL" region="15" clubid="1274" name="Kaliski Klub Sportowy  ,,Włókniarz&apos;&apos; 1925 Kalisz">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Szymański" birthdate="2005-05-06" gender="M" nation="POL" license="105415700007" swrid="4945641" athleteid="1275">
              <RESULTS>
                <RESULT eventid="1075" points="480" reactiontime="+80" swimtime="00:00:26.70" resultid="1276" heatid="2969" lane="6" entrytime="00:00:26.90" entrycourse="LCM" />
                <RESULT eventid="1091" points="409" reactiontime="+76" swimtime="00:01:06.65" resultid="1277" heatid="2981" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="553" reactiontime="+76" swimtime="00:02:16.30" resultid="1278" heatid="3028" lane="4" entrytime="00:02:17.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:06.52" />
                    <SPLIT distance="150" swimtime="00:01:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="549" reactiontime="+68" swimtime="00:01:03.30" resultid="1279" heatid="3065" lane="6" entrytime="00:01:03.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="KS Warszawianka" version="11.49155">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" phone="+41 99 999 99 99" fax="+41 99 999 99 99" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Warszawa" name="Letnie Mistrzostwa Polski w pływaniu Masters" course="LCM" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2017-06-16" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Warszawa" nation="POL" />
      <POINTTABLE pointtableid="3010" name="FINA Point Scoring" version="2017" />
      <SESSIONS>
        <SESSION date="2017-06-16" daytime="10:00" endtime="15:12" name="I Blok" number="1" warmupfrom="09:00" warmupuntil="09:50">
          <EVENTS>
            <EVENT eventid="1059" daytime="10:00" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1738" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3191" />
                    <RANKING order="2" place="-1" resultid="10122" />
                    <RANKING order="3" place="-1" resultid="10553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1739" agemax="29" agemin="25" name="Kat A - 25-29" />
                <AGEGROUP agegroupid="1740" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9866" />
                    <RANKING order="2" place="2" resultid="6442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1741" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3862" />
                    <RANKING order="2" place="2" resultid="7573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1742" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7901" />
                    <RANKING order="2" place="2" resultid="9358" />
                    <RANKING order="3" place="3" resultid="7652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1743" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8788" />
                    <RANKING order="2" place="2" resultid="7565" />
                    <RANKING order="3" place="-1" resultid="3235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1744" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1745" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6661" />
                    <RANKING order="2" place="2" resultid="6447" />
                    <RANKING order="3" place="3" resultid="9592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1746" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6680" />
                    <RANKING order="2" place="2" resultid="3201" />
                    <RANKING order="3" place="3" resultid="9602" />
                    <RANKING order="4" place="4" resultid="7561" />
                    <RANKING order="5" place="5" resultid="6454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1747" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4576" />
                    <RANKING order="2" place="2" resultid="8569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1748" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1749" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="1750" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="1752" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="1753" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="1751" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10665" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10666" daytime="10:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10667" daytime="10:42" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1128" daytime="13:16" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2331" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="10303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2332" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7061" />
                    <RANKING order="2" place="2" resultid="6848" />
                    <RANKING order="3" place="3" resultid="8219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2333" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8368" />
                    <RANKING order="2" place="2" resultid="6954" />
                    <RANKING order="3" place="3" resultid="10946" />
                    <RANKING order="4" place="4" resultid="7610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2334" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8573" />
                    <RANKING order="2" place="2" resultid="3187" />
                    <RANKING order="3" place="3" resultid="6886" />
                    <RANKING order="4" place="4" resultid="10640" />
                    <RANKING order="5" place="5" resultid="9372" />
                    <RANKING order="6" place="6" resultid="8361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2335" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6635" />
                    <RANKING order="2" place="2" resultid="6400" />
                    <RANKING order="3" place="3" resultid="6571" />
                    <RANKING order="4" place="4" resultid="9513" />
                    <RANKING order="5" place="5" resultid="6908" />
                    <RANKING order="6" place="6" resultid="8052" />
                    <RANKING order="7" place="7" resultid="10277" />
                    <RANKING order="8" place="8" resultid="8238" />
                    <RANKING order="9" place="9" resultid="10110" />
                    <RANKING order="10" place="10" resultid="7668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2336" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7409" />
                    <RANKING order="2" place="2" resultid="10079" />
                    <RANKING order="3" place="3" resultid="9783" />
                    <RANKING order="4" place="4" resultid="7622" />
                    <RANKING order="5" place="5" resultid="9420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2337" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6523" />
                    <RANKING order="2" place="2" resultid="7402" />
                    <RANKING order="3" place="3" resultid="8536" />
                    <RANKING order="4" place="4" resultid="7605" />
                    <RANKING order="5" place="5" resultid="9446" />
                    <RANKING order="6" place="6" resultid="7533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2338" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9115" />
                    <RANKING order="2" place="2" resultid="8044" />
                    <RANKING order="3" place="3" resultid="6758" />
                    <RANKING order="4" place="4" resultid="6403" />
                    <RANKING order="5" place="5" resultid="7394" />
                    <RANKING order="6" place="6" resultid="7940" />
                    <RANKING order="7" place="-1" resultid="7575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2339" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10265" />
                    <RANKING order="2" place="2" resultid="9542" />
                    <RANKING order="3" place="3" resultid="9803" />
                    <RANKING order="4" place="4" resultid="8093" />
                    <RANKING order="5" place="-1" resultid="9516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2340" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2341" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2342" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2343" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2344" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2345" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2346" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10675" daytime="13:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10676" daytime="14:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10677" daytime="14:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10678" daytime="14:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10679" daytime="15:18" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1098" daytime="10:58" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2299" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10302" />
                    <RANKING order="2" place="2" resultid="3622" />
                    <RANKING order="3" place="3" resultid="6472" />
                    <RANKING order="4" place="-1" resultid="10112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2300" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3640" />
                    <RANKING order="2" place="2" resultid="7767" />
                    <RANKING order="3" place="3" resultid="3837" />
                    <RANKING order="4" place="4" resultid="7738" />
                    <RANKING order="5" place="5" resultid="7068" />
                    <RANKING order="6" place="6" resultid="3517" />
                    <RANKING order="7" place="-1" resultid="10564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2301" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9102" />
                    <RANKING order="2" place="2" resultid="8832" />
                    <RANKING order="3" place="3" resultid="7152" />
                    <RANKING order="4" place="4" resultid="8587" />
                    <RANKING order="5" place="5" resultid="6054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2302" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9583" />
                    <RANKING order="2" place="2" resultid="8440" />
                    <RANKING order="3" place="3" resultid="7637" />
                    <RANKING order="4" place="4" resultid="8974" />
                    <RANKING order="5" place="5" resultid="8327" />
                    <RANKING order="6" place="6" resultid="8337" />
                    <RANKING order="7" place="7" resultid="6910" />
                    <RANKING order="8" place="-1" resultid="10287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2303" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7642" />
                    <RANKING order="2" place="2" resultid="9095" />
                    <RANKING order="3" place="3" resultid="8005" />
                    <RANKING order="4" place="4" resultid="8246" />
                    <RANKING order="5" place="-1" resultid="3853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2304" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8644" />
                    <RANKING order="2" place="2" resultid="3291" />
                    <RANKING order="3" place="3" resultid="8296" />
                    <RANKING order="4" place="4" resultid="8225" />
                    <RANKING order="5" place="5" resultid="6738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2305" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7581" />
                    <RANKING order="2" place="2" resultid="7395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2306" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9340" />
                    <RANKING order="2" place="2" resultid="7615" />
                    <RANKING order="3" place="3" resultid="8510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2307" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8980" />
                    <RANKING order="2" place="2" resultid="4558" />
                    <RANKING order="3" place="3" resultid="7993" />
                    <RANKING order="4" place="4" resultid="6378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2308" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8331" />
                    <RANKING order="2" place="2" resultid="8060" />
                    <RANKING order="3" place="3" resultid="8945" />
                    <RANKING order="4" place="4" resultid="9029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2309" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7771" />
                    <RANKING order="2" place="2" resultid="8577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2310" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6642" />
                    <RANKING order="2" place="-1" resultid="7970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2311" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2312" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2313" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2314" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10668" daytime="10:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10669" daytime="11:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10670" daytime="11:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10671" daytime="12:09" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10672" daytime="12:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10673" daytime="12:34" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="12:45" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2315" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2316" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7756" />
                    <RANKING order="2" place="2" resultid="3507" />
                    <RANKING order="3" place="-1" resultid="3630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2317" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9857" />
                    <RANKING order="2" place="2" resultid="9344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2318" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2319" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2320" agemax="49" agemin="45" name="Kat E 45-49" />
                <AGEGROUP agegroupid="2321" agemax="54" agemin="50" name="Kat F 50-54" />
                <AGEGROUP agegroupid="2322" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2323" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2324" agemax="69" agemin="65" name="Kat I 65-69" />
                <AGEGROUP agegroupid="2325" agemax="74" agemin="70" name="Kat J 70-74" />
                <AGEGROUP agegroupid="2326" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2327" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2328" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2329" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2330" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10674" daytime="12:45" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2017-06-16" daytime="16:00" endtime="19:14" name="II Blok" number="2" warmupfrom="14:30" warmupuntil="15:45">
          <EVENTS>
            <EVENT eventid="1160" daytime="16:12" gender="M" number="6" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2363" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7081" />
                    <RANKING order="2" place="2" resultid="8415" />
                    <RANKING order="3" place="3" resultid="6845" />
                    <RANKING order="4" place="4" resultid="10311" />
                    <RANKING order="5" place="5" resultid="10954" />
                    <RANKING order="6" place="6" resultid="10644" />
                    <RANKING order="7" place="7" resultid="7596" />
                    <RANKING order="8" place="8" resultid="6473" />
                    <RANKING order="9" place="9" resultid="10262" />
                    <RANKING order="10" place="10" resultid="9828" />
                    <RANKING order="11" place="11" resultid="10230" />
                    <RANKING order="12" place="12" resultid="3850" />
                    <RANKING order="13" place="-1" resultid="10113" />
                    <RANKING order="14" place="-1" resultid="10304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2364" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6330" />
                    <RANKING order="2" place="2" resultid="7590" />
                    <RANKING order="3" place="3" resultid="7008" />
                    <RANKING order="4" place="4" resultid="10292" />
                    <RANKING order="5" place="5" resultid="6813" />
                    <RANKING order="6" place="6" resultid="7739" />
                    <RANKING order="7" place="7" resultid="6296" />
                    <RANKING order="8" place="8" resultid="8468" />
                    <RANKING order="9" place="9" resultid="7089" />
                    <RANKING order="10" place="10" resultid="6859" />
                    <RANKING order="11" place="11" resultid="3518" />
                    <RANKING order="12" place="12" resultid="3838" />
                    <RANKING order="13" place="13" resultid="7136" />
                    <RANKING order="14" place="14" resultid="9399" />
                    <RANKING order="15" place="15" resultid="6919" />
                    <RANKING order="16" place="16" resultid="7131" />
                    <RANKING order="17" place="17" resultid="9416" />
                    <RANKING order="18" place="-1" resultid="6854" />
                    <RANKING order="19" place="-1" resultid="7012" />
                    <RANKING order="20" place="-1" resultid="7141" />
                    <RANKING order="21" place="-1" resultid="8220" />
                    <RANKING order="22" place="-1" resultid="9909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2365" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6798" />
                    <RANKING order="2" place="2" resultid="6796" />
                    <RANKING order="3" place="3" resultid="9224" />
                    <RANKING order="4" place="4" resultid="7908" />
                    <RANKING order="5" place="5" resultid="8967" />
                    <RANKING order="6" place="6" resultid="3875" />
                    <RANKING order="7" place="7" resultid="6800" />
                    <RANKING order="8" place="8" resultid="9875" />
                    <RANKING order="9" place="9" resultid="6881" />
                    <RANKING order="10" place="10" resultid="9806" />
                    <RANKING order="11" place="11" resultid="9889" />
                    <RANKING order="12" place="12" resultid="8552" />
                    <RANKING order="13" place="13" resultid="6810" />
                    <RANKING order="14" place="14" resultid="7790" />
                    <RANKING order="15" place="15" resultid="6902" />
                    <RANKING order="16" place="16" resultid="7092" />
                    <RANKING order="17" place="17" resultid="3826" />
                    <RANKING order="18" place="18" resultid="6955" />
                    <RANKING order="19" place="19" resultid="8856" />
                    <RANKING order="20" place="20" resultid="6302" />
                    <RANKING order="21" place="21" resultid="10947" />
                    <RANKING order="22" place="22" resultid="7611" />
                    <RANKING order="23" place="23" resultid="8602" />
                    <RANKING order="24" place="24" resultid="3890" />
                    <RANKING order="25" place="25" resultid="10568" />
                    <RANKING order="26" place="26" resultid="9818" />
                    <RANKING order="27" place="-1" resultid="8455" />
                    <RANKING order="28" place="-1" resultid="9442" />
                    <RANKING order="29" place="-1" resultid="9795" />
                    <RANKING order="30" place="-1" resultid="9897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2366" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8651" />
                    <RANKING order="2" place="2" resultid="9529" />
                    <RANKING order="3" place="3" resultid="6658" />
                    <RANKING order="4" place="4" resultid="6395" />
                    <RANKING order="5" place="5" resultid="9880" />
                    <RANKING order="6" place="6" resultid="8904" />
                    <RANKING order="7" place="7" resultid="8441" />
                    <RANKING order="8" place="8" resultid="9433" />
                    <RANKING order="9" place="9" resultid="6868" />
                    <RANKING order="10" place="10" resultid="6898" />
                    <RANKING order="11" place="11" resultid="6519" />
                    <RANKING order="12" place="12" resultid="3188" />
                    <RANKING order="13" place="13" resultid="6809" />
                    <RANKING order="14" place="14" resultid="9611" />
                    <RANKING order="15" place="15" resultid="6873" />
                    <RANKING order="16" place="16" resultid="9395" />
                    <RANKING order="17" place="17" resultid="7638" />
                    <RANKING order="18" place="18" resultid="8559" />
                    <RANKING order="19" place="19" resultid="8525" />
                    <RANKING order="20" place="20" resultid="6911" />
                    <RANKING order="21" place="21" resultid="7000" />
                    <RANKING order="22" place="22" resultid="7650" />
                    <RANKING order="23" place="23" resultid="10039" />
                    <RANKING order="24" place="24" resultid="6997" />
                    <RANKING order="25" place="25" resultid="7018" />
                    <RANKING order="26" place="26" resultid="8606" />
                    <RANKING order="27" place="27" resultid="3271" />
                    <RANKING order="28" place="28" resultid="10659" />
                    <RANKING order="29" place="-1" resultid="7020" />
                    <RANKING order="30" place="-1" resultid="8975" />
                    <RANKING order="31" place="-1" resultid="9456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2367" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6776" />
                    <RANKING order="2" place="2" resultid="8006" />
                    <RANKING order="3" place="3" resultid="7643" />
                    <RANKING order="4" place="4" resultid="8076" />
                    <RANKING order="5" place="5" resultid="8257" />
                    <RANKING order="6" place="6" resultid="6811" />
                    <RANKING order="7" place="7" resultid="10236" />
                    <RANKING order="8" place="8" resultid="9381" />
                    <RANKING order="9" place="9" resultid="6576" />
                    <RANKING order="10" place="10" resultid="8016" />
                    <RANKING order="11" place="11" resultid="6651" />
                    <RANKING order="12" place="12" resultid="8247" />
                    <RANKING order="13" place="13" resultid="8448" />
                    <RANKING order="14" place="14" resultid="8011" />
                    <RANKING order="15" place="14" resultid="8617" />
                    <RANKING order="16" place="16" resultid="8593" />
                    <RANKING order="17" place="17" resultid="8487" />
                    <RANKING order="18" place="18" resultid="3854" />
                    <RANKING order="19" place="19" resultid="8239" />
                    <RANKING order="20" place="20" resultid="6909" />
                    <RANKING order="21" place="21" resultid="10252" />
                    <RANKING order="22" place="22" resultid="8462" />
                    <RANKING order="23" place="23" resultid="7669" />
                    <RANKING order="24" place="24" resultid="9791" />
                    <RANKING order="25" place="-1" resultid="6966" />
                    <RANKING order="26" place="-1" resultid="6968" />
                    <RANKING order="27" place="-1" resultid="7794" />
                    <RANKING order="28" place="-1" resultid="8465" />
                    <RANKING order="29" place="-1" resultid="10157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2368" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6978" />
                    <RANKING order="2" place="2" resultid="8539" />
                    <RANKING order="3" place="3" resultid="6983" />
                    <RANKING order="4" place="4" resultid="8645" />
                    <RANKING order="5" place="5" resultid="10167" />
                    <RANKING order="6" place="6" resultid="4567" />
                    <RANKING order="7" place="7" resultid="3292" />
                    <RANKING order="8" place="8" resultid="7414" />
                    <RANKING order="9" place="9" resultid="8198" />
                    <RANKING order="10" place="10" resultid="10080" />
                    <RANKING order="11" place="11" resultid="8251" />
                    <RANKING order="12" place="12" resultid="8226" />
                    <RANKING order="13" place="13" resultid="8424" />
                    <RANKING order="14" place="14" resultid="7021" />
                    <RANKING order="15" place="15" resultid="8216" />
                    <RANKING order="16" place="15" resultid="10654" />
                    <RANKING order="17" place="17" resultid="8474" />
                    <RANKING order="18" place="18" resultid="9421" />
                    <RANKING order="19" place="19" resultid="9813" />
                    <RANKING order="20" place="20" resultid="3886" />
                    <RANKING order="21" place="21" resultid="9404" />
                    <RANKING order="22" place="-1" resultid="3301" />
                    <RANKING order="23" place="-1" resultid="7410" />
                    <RANKING order="24" place="-1" resultid="8614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2369" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6282" />
                    <RANKING order="2" place="2" resultid="6434" />
                    <RANKING order="3" place="3" resultid="8518" />
                    <RANKING order="4" place="4" resultid="10576" />
                    <RANKING order="5" place="5" resultid="6427" />
                    <RANKING order="6" place="6" resultid="6524" />
                    <RANKING order="7" place="7" resultid="6534" />
                    <RANKING order="8" place="8" resultid="8597" />
                    <RANKING order="9" place="9" resultid="6806" />
                    <RANKING order="10" place="10" resultid="7582" />
                    <RANKING order="11" place="11" resultid="7396" />
                    <RANKING order="12" place="12" resultid="9447" />
                    <RANKING order="13" place="13" resultid="7403" />
                    <RANKING order="14" place="14" resultid="6630" />
                    <RANKING order="15" place="15" resultid="7606" />
                    <RANKING order="16" place="16" resultid="6328" />
                    <RANKING order="17" place="17" resultid="7534" />
                    <RANKING order="18" place="17" resultid="8497" />
                    <RANKING order="19" place="19" resultid="10281" />
                    <RANKING order="20" place="20" resultid="9787" />
                    <RANKING order="21" place="21" resultid="9808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2370" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8503" />
                    <RANKING order="2" place="2" resultid="9916" />
                    <RANKING order="3" place="3" resultid="9619" />
                    <RANKING order="4" place="4" resultid="6689" />
                    <RANKING order="5" place="5" resultid="7633" />
                    <RANKING order="6" place="6" resultid="9116" />
                    <RANKING order="7" place="7" resultid="8775" />
                    <RANKING order="8" place="8" resultid="8950" />
                    <RANKING order="9" place="9" resultid="7390" />
                    <RANKING order="10" place="10" resultid="6759" />
                    <RANKING order="11" place="11" resultid="6349" />
                    <RANKING order="12" place="12" resultid="8511" />
                    <RANKING order="13" place="-1" resultid="9378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2371" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10329" />
                    <RANKING order="2" place="2" resultid="9926" />
                    <RANKING order="3" place="3" resultid="8981" />
                    <RANKING order="4" place="4" resultid="10266" />
                    <RANKING order="5" place="5" resultid="6771" />
                    <RANKING order="6" place="6" resultid="6379" />
                    <RANKING order="7" place="7" resultid="7382" />
                    <RANKING order="8" place="8" resultid="6788" />
                    <RANKING order="9" place="9" resultid="7525" />
                    <RANKING order="10" place="10" resultid="6502" />
                    <RANKING order="11" place="11" resultid="7105" />
                    <RANKING order="12" place="12" resultid="8895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2372" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8332" />
                    <RANKING order="2" place="2" resultid="8061" />
                    <RANKING order="3" place="3" resultid="8781" />
                    <RANKING order="4" place="4" resultid="9055" />
                    <RANKING order="5" place="5" resultid="7378" />
                    <RANKING order="6" place="6" resultid="8785" />
                    <RANKING order="7" place="7" resultid="9030" />
                    <RANKING order="8" place="-1" resultid="6527" />
                    <RANKING order="9" place="-1" resultid="7551" />
                    <RANKING order="10" place="-1" resultid="7911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2373" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8922" />
                    <RANKING order="2" place="2" resultid="7772" />
                    <RANKING order="3" place="3" resultid="7477" />
                    <RANKING order="4" place="4" resultid="6614" />
                    <RANKING order="5" place="5" resultid="7374" />
                    <RANKING order="6" place="6" resultid="8578" />
                    <RANKING order="7" place="7" resultid="7985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2374" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8209" />
                    <RANKING order="2" place="2" resultid="9060" />
                    <RANKING order="3" place="3" resultid="8431" />
                    <RANKING order="4" place="4" resultid="8345" />
                    <RANKING order="5" place="5" resultid="6643" />
                    <RANKING order="6" place="-1" resultid="7971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2375" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7749" />
                    <RANKING order="2" place="2" resultid="8350" />
                    <RANKING order="3" place="3" resultid="11055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2376" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3242" />
                    <RANKING order="2" place="2" resultid="3159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2377" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2378" agemax="99" agemin="95" name="Kat O 95-99">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8881" />
                    <RANKING order="2" place="-1" resultid="7322" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10689" daytime="16:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10690" daytime="16:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10691" daytime="16:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10692" daytime="16:17" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10693" daytime="16:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10694" daytime="16:19" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10695" daytime="16:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10696" daytime="16:21" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10697" daytime="16:22" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10698" daytime="16:23" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10699" daytime="16:24" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10700" daytime="16:25" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="10701" daytime="16:26" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="10702" daytime="16:27" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="10703" daytime="16:28" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="10704" daytime="16:29" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="10705" daytime="16:30" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="10706" daytime="16:31" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="10707" daytime="16:32" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="10708" daytime="16:33" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="10709" daytime="16:34" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="10710" daytime="16:35" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="10711" daytime="16:36" number="23" order="23" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1175" daytime="16:37" gender="F" number="7" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2379" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9495" />
                    <RANKING order="2" place="2" resultid="7946" />
                    <RANKING order="3" place="3" resultid="3831" />
                    <RANKING order="4" place="4" resultid="7677" />
                    <RANKING order="5" place="5" resultid="7663" />
                    <RANKING order="6" place="6" resultid="3193" />
                    <RANKING order="7" place="-1" resultid="10124" />
                    <RANKING order="8" place="-1" resultid="10554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2380" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3222" />
                    <RANKING order="2" place="2" resultid="7026" />
                    <RANKING order="3" place="3" resultid="7758" />
                    <RANKING order="4" place="4" resultid="3509" />
                    <RANKING order="5" place="-1" resultid="3631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2381" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6782" />
                    <RANKING order="2" place="2" resultid="8374" />
                    <RANKING order="3" place="3" resultid="6590" />
                    <RANKING order="4" place="4" resultid="9858" />
                    <RANKING order="5" place="5" resultid="9498" />
                    <RANKING order="6" place="6" resultid="10294" />
                    <RANKING order="7" place="7" resultid="8661" />
                    <RANKING order="8" place="8" resultid="9345" />
                    <RANKING order="9" place="9" resultid="10319" />
                    <RANKING order="10" place="10" resultid="9868" />
                    <RANKING order="11" place="11" resultid="8482" />
                    <RANKING order="12" place="-1" resultid="8547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2382" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7962" />
                    <RANKING order="2" place="2" resultid="3864" />
                    <RANKING order="3" place="3" resultid="6321" />
                    <RANKING order="4" place="4" resultid="8265" />
                    <RANKING order="5" place="5" resultid="10086" />
                    <RANKING order="6" place="6" resultid="8849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2383" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8954" />
                    <RANKING order="2" place="2" resultid="8827" />
                    <RANKING order="3" place="3" resultid="9805" />
                    <RANKING order="4" place="4" resultid="3284" />
                    <RANKING order="5" place="5" resultid="6765" />
                    <RANKING order="6" place="6" resultid="6654" />
                    <RANKING order="7" place="7" resultid="9823" />
                    <RANKING order="8" place="-1" resultid="6988" />
                    <RANKING order="9" place="-1" resultid="7654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2384" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7354" />
                    <RANKING order="2" place="2" resultid="8959" />
                    <RANKING order="3" place="3" resultid="3646" />
                    <RANKING order="4" place="4" resultid="8621" />
                    <RANKING order="5" place="5" resultid="6675" />
                    <RANKING order="6" place="6" resultid="6638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2385" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6648" />
                    <RANKING order="2" place="2" resultid="8070" />
                    <RANKING order="3" place="3" resultid="6356" />
                    <RANKING order="4" place="4" resultid="6288" />
                    <RANKING order="5" place="-1" resultid="6410" />
                    <RANKING order="6" place="-1" resultid="3793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2386" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8938" />
                    <RANKING order="2" place="2" resultid="8087" />
                    <RANKING order="3" place="3" resultid="6663" />
                    <RANKING order="4" place="4" resultid="9351" />
                    <RANKING order="5" place="5" resultid="9594" />
                    <RANKING order="6" place="6" resultid="6448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2387" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9578" />
                    <RANKING order="2" place="2" resultid="7340" />
                    <RANKING order="3" place="3" resultid="10093" />
                    <RANKING order="4" place="4" resultid="6682" />
                    <RANKING order="5" place="5" resultid="3202" />
                    <RANKING order="6" place="-1" resultid="3213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2388" agemax="69" agemin="65" name="Kat I 65-69" />
                <AGEGROUP agegroupid="2389" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2390" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2391" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2392" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2393" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2394" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10712" daytime="16:37" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10713" daytime="16:43" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10714" daytime="16:49" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10715" daytime="16:53" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10716" daytime="16:57" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10717" daytime="17:00" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10718" daytime="17:04" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1144" daytime="16:00" gender="F" number="5" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2347" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7945" />
                    <RANKING order="2" place="2" resultid="9494" />
                    <RANKING order="3" place="3" resultid="3821" />
                    <RANKING order="4" place="4" resultid="10298" />
                    <RANKING order="5" place="5" resultid="9374" />
                    <RANKING order="6" place="6" resultid="3307" />
                    <RANKING order="7" place="7" resultid="3192" />
                    <RANKING order="8" place="8" resultid="9438" />
                    <RANKING order="9" place="-1" resultid="10123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2348" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3221" />
                    <RANKING order="2" place="2" resultid="8636" />
                    <RANKING order="3" place="3" resultid="7757" />
                    <RANKING order="4" place="4" resultid="3508" />
                    <RANKING order="5" place="5" resultid="11060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2349" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7369" />
                    <RANKING order="2" place="2" resultid="6781" />
                    <RANKING order="3" place="3" resultid="8373" />
                    <RANKING order="4" place="4" resultid="9844" />
                    <RANKING order="5" place="5" resultid="8610" />
                    <RANKING order="6" place="6" resultid="7078" />
                    <RANKING order="7" place="7" resultid="8913" />
                    <RANKING order="8" place="8" resultid="9867" />
                    <RANKING order="9" place="9" resultid="9849" />
                    <RANKING order="10" place="10" resultid="10318" />
                    <RANKING order="11" place="11" resultid="3845" />
                    <RANKING order="12" place="12" resultid="7004" />
                    <RANKING order="13" place="13" resultid="6443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2350" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7961" />
                    <RANKING order="2" place="2" resultid="6320" />
                    <RANKING order="3" place="3" resultid="6880" />
                    <RANKING order="4" place="4" resultid="3863" />
                    <RANKING order="5" place="5" resultid="7365" />
                    <RANKING order="6" place="6" resultid="8264" />
                    <RANKING order="7" place="7" resultid="7659" />
                    <RANKING order="8" place="8" resultid="9390" />
                    <RANKING order="9" place="9" resultid="9423" />
                    <RANKING order="10" place="10" resultid="8848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2351" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6315" />
                    <RANKING order="2" place="2" resultid="9487" />
                    <RANKING order="3" place="3" resultid="8291" />
                    <RANKING order="4" place="4" resultid="6581" />
                    <RANKING order="5" place="5" resultid="6586" />
                    <RANKING order="6" place="6" resultid="7653" />
                    <RANKING order="7" place="7" resultid="9804" />
                    <RANKING order="8" place="8" resultid="9411" />
                    <RANKING order="9" place="9" resultid="3257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2352" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6670" />
                    <RANKING order="2" place="2" resultid="10103" />
                    <RANKING order="3" place="3" resultid="6674" />
                    <RANKING order="4" place="4" resultid="8620" />
                    <RANKING order="5" place="5" resultid="6637" />
                    <RANKING order="6" place="6" resultid="7566" />
                    <RANKING order="7" place="-1" resultid="3236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2353" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6604" />
                    <RANKING order="2" place="2" resultid="6355" />
                    <RANKING order="3" place="3" resultid="10652" />
                    <RANKING order="4" place="4" resultid="8069" />
                    <RANKING order="5" place="5" resultid="6409" />
                    <RANKING order="6" place="-1" resultid="3792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2354" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8937" />
                    <RANKING order="2" place="2" resultid="8929" />
                    <RANKING order="3" place="3" resultid="6662" />
                    <RANKING order="4" place="4" resultid="7350" />
                    <RANKING order="5" place="5" resultid="6482" />
                    <RANKING order="6" place="6" resultid="9593" />
                    <RANKING order="7" place="7" resultid="6489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2355" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7334" />
                    <RANKING order="2" place="2" resultid="6681" />
                    <RANKING order="3" place="3" resultid="3212" />
                    <RANKING order="4" place="4" resultid="9603" />
                    <RANKING order="5" place="5" resultid="10605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2356" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4577" />
                    <RANKING order="2" place="2" resultid="8771" />
                    <RANKING order="3" place="3" resultid="7481" />
                    <RANKING order="4" place="4" resultid="9068" />
                    <RANKING order="5" place="5" resultid="8570" />
                    <RANKING order="6" place="6" resultid="3651" />
                    <RANKING order="7" place="-1" resultid="7326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2357" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8768" />
                    <RANKING order="2" place="2" resultid="6622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2358" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2359" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2360" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2361" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2362" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10680" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10681" daytime="16:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10682" daytime="16:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10683" daytime="16:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10684" daytime="16:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10685" daytime="16:07" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10686" daytime="16:08" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10687" daytime="16:09" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10688" daytime="16:11" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="17:53" number="9" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1220" agemax="119" agemin="100" name="Kat A 100-119">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="159" agemin="120" name="Kat B 120-159">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8665" />
                    <RANKING order="2" place="2" resultid="6922" />
                    <RANKING order="3" place="3" resultid="9905" />
                    <RANKING order="4" place="4" resultid="3894" />
                    <RANKING order="5" place="5" resultid="7685" />
                    <RANKING order="6" place="6" resultid="8864" />
                    <RANKING order="7" place="7" resultid="9457" />
                    <RANKING order="8" place="-1" resultid="9458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="199" agemin="160" name="Kat C 160-199">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6696" />
                    <RANKING order="2" place="2" resultid="7427" />
                    <RANKING order="3" place="3" resultid="9002" />
                    <RANKING order="4" place="4" resultid="8666" />
                    <RANKING order="5" place="5" resultid="8667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="239" agemin="200" name="Kat D 200-239">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7425" />
                    <RANKING order="2" place="2" resultid="6698" />
                    <RANKING order="3" place="3" resultid="9641" />
                    <RANKING order="4" place="4" resultid="6514" />
                    <RANKING order="5" place="5" resultid="3313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="279" agemin="240" name="Kat E 240-279">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9003" />
                    <RANKING order="2" place="2" resultid="7423" />
                    <RANKING order="3" place="3" resultid="8799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="-1" agemin="280" name="Kat F 280 +">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8798" />
                    <RANKING order="2" place="-1" resultid="9907" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10731" daytime="17:53" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10732" daytime="17:57" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10733" daytime="18:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1190" daytime="17:08" gender="M" number="8" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2395" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9518" />
                    <RANKING order="2" place="2" resultid="7082" />
                    <RANKING order="3" place="3" resultid="3623" />
                    <RANKING order="4" place="4" resultid="10645" />
                    <RANKING order="5" place="5" resultid="6474" />
                    <RANKING order="6" place="6" resultid="9829" />
                    <RANKING order="7" place="-1" resultid="10114" />
                    <RANKING order="8" place="-1" resultid="10305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2396" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7768" />
                    <RANKING order="2" place="2" resultid="7069" />
                    <RANKING order="3" place="3" resultid="7601" />
                    <RANKING order="4" place="4" resultid="3641" />
                    <RANKING order="5" place="5" resultid="7062" />
                    <RANKING order="6" place="6" resultid="6849" />
                    <RANKING order="7" place="7" resultid="3519" />
                    <RANKING order="8" place="8" resultid="6860" />
                    <RANKING order="9" place="-1" resultid="6855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2397" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6801" />
                    <RANKING order="2" place="2" resultid="8833" />
                    <RANKING order="3" place="3" resultid="6892" />
                    <RANKING order="4" place="4" resultid="3876" />
                    <RANKING order="5" place="5" resultid="6903" />
                    <RANKING order="6" place="6" resultid="9890" />
                    <RANKING order="7" place="7" resultid="8588" />
                    <RANKING order="8" place="8" resultid="7626" />
                    <RANKING order="9" place="9" resultid="8857" />
                    <RANKING order="10" place="-1" resultid="9796" />
                    <RANKING order="11" place="-1" resultid="6956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2398" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9584" />
                    <RANKING order="2" place="2" resultid="9881" />
                    <RANKING order="3" place="3" resultid="8905" />
                    <RANKING order="4" place="4" resultid="6887" />
                    <RANKING order="5" place="5" resultid="8841" />
                    <RANKING order="6" place="6" resultid="9427" />
                    <RANKING order="7" place="7" resultid="9434" />
                    <RANKING order="8" place="8" resultid="6508" />
                    <RANKING order="9" place="9" resultid="8338" />
                    <RANKING order="10" place="10" resultid="6912" />
                    <RANKING order="11" place="11" resultid="8362" />
                    <RANKING order="12" place="12" resultid="3272" />
                    <RANKING order="13" place="-1" resultid="7001" />
                    <RANKING order="14" place="-1" resultid="9612" />
                    <RANKING order="15" place="-1" resultid="10288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2399" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8077" />
                    <RANKING order="2" place="2" resultid="7644" />
                    <RANKING order="3" place="3" resultid="8258" />
                    <RANKING order="4" place="4" resultid="8449" />
                    <RANKING order="5" place="5" resultid="10237" />
                    <RANKING order="6" place="6" resultid="9922" />
                    <RANKING order="7" place="7" resultid="7156" />
                    <RANKING order="8" place="8" resultid="8021" />
                    <RANKING order="9" place="9" resultid="8563" />
                    <RANKING order="10" place="10" resultid="10278" />
                    <RANKING order="11" place="11" resultid="10253" />
                    <RANKING order="12" place="12" resultid="3855" />
                    <RANKING order="13" place="-1" resultid="8053" />
                    <RANKING order="14" place="-1" resultid="8488" />
                    <RANKING order="15" place="-1" resultid="10272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2400" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7781" />
                    <RANKING order="2" place="2" resultid="3787" />
                    <RANKING order="3" place="3" resultid="8232" />
                    <RANKING order="4" place="4" resultid="10081" />
                    <RANKING order="5" place="5" resultid="8227" />
                    <RANKING order="6" place="6" resultid="6739" />
                    <RANKING order="7" place="7" resultid="4568" />
                    <RANKING order="8" place="8" resultid="8475" />
                    <RANKING order="9" place="9" resultid="9405" />
                    <RANKING order="10" place="-1" resultid="3293" />
                    <RANKING order="11" place="-1" resultid="6420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2401" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6428" />
                    <RANKING order="2" place="2" resultid="10162" />
                    <RANKING order="3" place="3" resultid="8519" />
                    <RANKING order="4" place="4" resultid="6283" />
                    <RANKING order="5" place="5" resultid="10577" />
                    <RANKING order="6" place="6" resultid="7583" />
                    <RANKING order="7" place="7" resultid="7404" />
                    <RANKING order="8" place="8" resultid="8598" />
                    <RANKING order="9" place="9" resultid="9448" />
                    <RANKING order="10" place="10" resultid="6342" />
                    <RANKING order="11" place="11" resultid="10282" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2402" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8504" />
                    <RANKING order="2" place="2" resultid="7745" />
                    <RANKING order="3" place="3" resultid="9341" />
                    <RANKING order="4" place="4" resultid="10616" />
                    <RANKING order="5" place="5" resultid="9624" />
                    <RANKING order="6" place="6" resultid="8045" />
                    <RANKING order="7" place="7" resultid="6404" />
                    <RANKING order="8" place="8" resultid="7941" />
                    <RANKING order="9" place="-1" resultid="6760" />
                    <RANKING order="10" place="-1" resultid="7545" />
                    <RANKING order="11" place="-1" resultid="7576" />
                    <RANKING order="12" place="-1" resultid="7616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2403" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10571" />
                    <RANKING order="2" place="2" resultid="8531" />
                    <RANKING order="3" place="3" resultid="7922" />
                    <RANKING order="4" place="4" resultid="6305" />
                    <RANKING order="5" place="5" resultid="7383" />
                    <RANKING order="6" place="6" resultid="4559" />
                    <RANKING order="7" place="7" resultid="8556" />
                    <RANKING order="8" place="8" resultid="6789" />
                    <RANKING order="9" place="9" resultid="7994" />
                    <RANKING order="10" place="10" resultid="8896" />
                    <RANKING order="11" place="11" resultid="8886" />
                    <RANKING order="12" place="-1" resultid="8982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2404" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8631" />
                    <RANKING order="2" place="2" resultid="8062" />
                    <RANKING order="3" place="3" resultid="8890" />
                    <RANKING order="4" place="4" resultid="8380" />
                    <RANKING order="5" place="5" resultid="9031" />
                    <RANKING order="6" place="6" resultid="9836" />
                    <RANKING order="7" place="7" resultid="8354" />
                    <RANKING order="8" place="-1" resultid="8458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2405" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7773" />
                    <RANKING order="2" place="2" resultid="6615" />
                    <RANKING order="3" place="3" resultid="7986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2406" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9061" />
                    <RANKING order="2" place="2" resultid="7972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2407" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2408" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2409" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2410" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10719" daytime="17:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10720" daytime="17:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10721" daytime="17:19" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10722" daytime="17:23" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10723" daytime="17:27" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10724" daytime="17:31" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10725" daytime="17:34" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10726" daytime="17:37" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10727" daytime="17:41" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10728" daytime="17:44" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10729" daytime="17:47" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10730" daytime="17:50" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2017-06-17" daytime="09:00" endtime="12:48" name="Blok III" number="3" warmupfrom="07:30" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="1272" daytime="09:49" gender="M" number="13" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2459" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6387" />
                    <RANKING order="2" place="2" resultid="9519" />
                    <RANKING order="3" place="3" resultid="3625" />
                    <RANKING order="4" place="4" resultid="10116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2460" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6814" />
                    <RANKING order="2" place="2" resultid="7070" />
                    <RANKING order="3" place="3" resultid="8221" />
                    <RANKING order="4" place="4" resultid="6298" />
                    <RANKING order="5" place="5" resultid="3520" />
                    <RANKING order="6" place="6" resultid="7137" />
                    <RANKING order="7" place="-1" resultid="6856" />
                    <RANKING order="8" place="-1" resultid="10565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2461" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8603" />
                    <RANKING order="2" place="2" resultid="8369" />
                    <RANKING order="3" place="3" resultid="6904" />
                    <RANKING order="4" place="4" resultid="7627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2462" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9585" />
                    <RANKING order="2" place="2" resultid="8906" />
                    <RANKING order="3" place="3" resultid="8560" />
                    <RANKING order="4" place="4" resultid="6874" />
                    <RANKING order="5" place="5" resultid="9613" />
                    <RANKING order="6" place="6" resultid="6913" />
                    <RANKING order="7" place="7" resultid="10560" />
                    <RANKING order="8" place="8" resultid="3251" />
                    <RANKING order="9" place="-1" resultid="10289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2463" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8007" />
                    <RANKING order="2" place="2" resultid="8450" />
                    <RANKING order="3" place="3" resultid="6610" />
                    <RANKING order="4" place="4" resultid="10620" />
                    <RANKING order="5" place="5" resultid="10255" />
                    <RANKING order="6" place="6" resultid="8055" />
                    <RANKING order="7" place="7" resultid="3182" />
                    <RANKING order="8" place="-1" resultid="10158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2464" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6421" />
                    <RANKING order="2" place="2" resultid="8233" />
                    <RANKING order="3" place="3" resultid="3294" />
                    <RANKING order="4" place="4" resultid="8228" />
                    <RANKING order="5" place="5" resultid="6740" />
                    <RANKING order="6" place="6" resultid="7787" />
                    <RANKING order="7" place="7" resultid="8253" />
                    <RANKING order="8" place="8" resultid="8476" />
                    <RANKING order="9" place="-1" resultid="6973" />
                    <RANKING order="10" place="-1" resultid="8297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2465" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8599" />
                    <RANKING order="2" place="2" resultid="7397" />
                    <RANKING order="3" place="3" resultid="8498" />
                    <RANKING order="4" place="4" resultid="6343" />
                    <RANKING order="5" place="5" resultid="10283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2466" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6536" />
                    <RANKING order="2" place="2" resultid="9625" />
                    <RANKING order="3" place="-1" resultid="7546" />
                    <RANKING order="4" place="-1" resultid="7577" />
                    <RANKING order="5" place="-1" resultid="8919" />
                    <RANKING order="6" place="-1" resultid="9107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2467" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10572" />
                    <RANKING order="2" place="2" resultid="7923" />
                    <RANKING order="3" place="3" resultid="9073" />
                    <RANKING order="4" place="4" resultid="6306" />
                    <RANKING order="5" place="5" resultid="8557" />
                    <RANKING order="6" place="6" resultid="9125" />
                    <RANKING order="7" place="-1" resultid="8094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2468" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8632" />
                    <RANKING order="2" place="2" resultid="8946" />
                    <RANKING order="3" place="3" resultid="8891" />
                    <RANKING order="4" place="4" resultid="7379" />
                    <RANKING order="5" place="5" resultid="3230" />
                    <RANKING order="6" place="-1" resultid="7556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2469" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7830" />
                    <RANKING order="2" place="2" resultid="7478" />
                    <RANKING order="3" place="3" resultid="7774" />
                    <RANKING order="4" place="4" resultid="7987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2470" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8757" />
                    <RANKING order="2" place="2" resultid="6371" />
                    <RANKING order="3" place="3" resultid="9063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2471" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2472" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2473" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2474" agemax="99" agemin="95" name="Kat O 95-99">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7323" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10757" daytime="09:49" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10758" daytime="09:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10759" daytime="10:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10760" daytime="10:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10761" daytime="10:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10762" daytime="10:12" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10763" daytime="10:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10764" daytime="10:19" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1317" daytime="11:10" gender="F" number="16" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2507" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6390" />
                    <RANKING order="2" place="2" resultid="7678" />
                    <RANKING order="3" place="3" resultid="3195" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2508" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3511" />
                    <RANKING order="2" place="-1" resultid="3633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2509" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9499" />
                    <RANKING order="2" place="2" resultid="9860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2510" agemax="39" agemin="35" name="Kat C 35-39" />
                <AGEGROUP agegroupid="2511" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2512" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2513" agemax="54" agemin="50" name="Kat F 50-54" />
                <AGEGROUP agegroupid="2514" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8931" />
                    <RANKING order="2" place="2" resultid="6449" />
                    <RANKING order="3" place="3" resultid="9596" />
                    <RANKING order="4" place="-1" resultid="6491" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2515" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2516" agemax="69" agemin="65" name="Kat I 65-69" />
                <AGEGROUP agegroupid="2517" agemax="74" agemin="70" name="Kat J 70-74" />
                <AGEGROUP agegroupid="2518" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2519" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2520" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2521" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2522" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10789" daytime="11:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10790" daytime="11:15" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1368" daytime="11:55" gender="M" number="19" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1369" agemax="119" agemin="100" name="Kat A 100-119">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7027" />
                    <RANKING order="2" place="2" resultid="6818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1370" agemax="159" agemin="120" name="Kat B 120-159">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7681" />
                    <RANKING order="2" place="2" resultid="6923" />
                    <RANKING order="3" place="3" resultid="8670" />
                    <RANKING order="4" place="4" resultid="9460" />
                    <RANKING order="5" place="5" resultid="6924" />
                    <RANKING order="6" place="6" resultid="3897" />
                    <RANKING order="7" place="7" resultid="7029" />
                    <RANKING order="8" place="-1" resultid="7689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1371" agemax="199" agemin="160" name="Kat C 160-199">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9642" />
                    <RANKING order="2" place="2" resultid="8995" />
                    <RANKING order="3" place="3" resultid="8669" />
                    <RANKING order="4" place="4" resultid="8029" />
                    <RANKING order="5" place="5" resultid="8272" />
                    <RANKING order="6" place="6" resultid="6699" />
                    <RANKING order="7" place="7" resultid="8388" />
                    <RANKING order="8" place="8" resultid="3315" />
                    <RANKING order="9" place="-1" resultid="7800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1372" agemax="239" agemin="200" name="Kat D 200-239">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8668" />
                    <RANKING order="2" place="2" resultid="7683" />
                    <RANKING order="3" place="3" resultid="7434" />
                    <RANKING order="4" place="-1" resultid="7684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1373" agemax="279" agemin="240" name="Kat E 240-279">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7431" />
                    <RANKING order="2" place="2" resultid="8997" />
                    <RANKING order="3" place="3" resultid="6700" />
                    <RANKING order="4" place="4" resultid="3316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1374" agemax="-1" agemin="280" name="Kat F 280 +">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8801" />
                    <RANKING order="2" place="2" resultid="9081" />
                    <RANKING order="3" place="3" resultid="8386" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10799" daytime="11:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10800" daytime="11:59" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10801" daytime="12:03" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10802" daytime="12:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1257" daytime="09:24" gender="F" number="12" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2443" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9386" />
                    <RANKING order="2" place="2" resultid="10126" />
                    <RANKING order="3" place="3" resultid="3308" />
                    <RANKING order="4" place="4" resultid="3194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2444" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3223" />
                    <RANKING order="2" place="2" resultid="3510" />
                    <RANKING order="3" place="-1" resultid="3632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2445" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8375" />
                    <RANKING order="2" place="2" resultid="9859" />
                    <RANKING order="3" place="3" resultid="6591" />
                    <RANKING order="4" place="4" resultid="8611" />
                    <RANKING order="5" place="5" resultid="9869" />
                    <RANKING order="6" place="6" resultid="8483" />
                    <RANKING order="7" place="7" resultid="9850" />
                    <RANKING order="8" place="8" resultid="3872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2446" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8267" />
                    <RANKING order="2" place="2" resultid="6496" />
                    <RANKING order="3" place="3" resultid="8851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2447" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6316" />
                    <RANKING order="2" place="2" resultid="9533" />
                    <RANKING order="3" place="3" resultid="3285" />
                    <RANKING order="4" place="4" resultid="6766" />
                    <RANKING order="5" place="5" resultid="6655" />
                    <RANKING order="6" place="6" resultid="7833" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2448" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7356" />
                    <RANKING order="2" place="2" resultid="3647" />
                    <RANKING order="3" place="3" resultid="8789" />
                    <RANKING order="4" place="4" resultid="8622" />
                    <RANKING order="5" place="5" resultid="3265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2449" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2450" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8939" />
                    <RANKING order="2" place="2" resultid="9352" />
                    <RANKING order="3" place="3" resultid="9595" />
                    <RANKING order="4" place="4" resultid="6490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2451" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9579" />
                    <RANKING order="2" place="2" resultid="7335" />
                    <RANKING order="3" place="3" resultid="7347" />
                    <RANKING order="4" place="4" resultid="8310" />
                    <RANKING order="5" place="5" resultid="9605" />
                    <RANKING order="6" place="6" resultid="7562" />
                    <RANKING order="7" place="7" resultid="10607" />
                    <RANKING order="8" place="-1" resultid="6456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2452" agemax="69" agemin="65" name="Kat I 65-69" />
                <AGEGROUP agegroupid="2453" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8760" />
                    <RANKING order="2" place="2" resultid="6624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2454" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2455" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2456" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2457" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2458" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10752" daytime="09:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10753" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10754" daytime="09:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10755" daytime="09:41" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10756" daytime="09:45" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1347" daytime="11:47" gender="F" number="18" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1362" agemax="119" agemin="100" name="Kat A 100-119" />
                <AGEGROUP agegroupid="1363" agemax="159" agemin="120" name="Kat B 120-159">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9903" />
                    <RANKING order="2" place="2" resultid="8866" />
                    <RANKING order="3" place="3" resultid="8671" />
                    <RANKING order="4" place="-1" resultid="11200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1364" agemax="199" agemin="160" name="Kat C 160-199">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7430" />
                    <RANKING order="2" place="2" resultid="3314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1365" agemax="239" agemin="200" name="Kat D 200-239">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8999" />
                    <RANKING order="2" place="2" resultid="6701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1366" agemax="279" agemin="240" name="Kat E 240-279">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8800" />
                    <RANKING order="2" place="2" resultid="7429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1367" agemax="-1" agemin="280" name="Kat F 280 +" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10797" daytime="11:47" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10798" daytime="11:51" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1287" daytime="10:22" gender="F" number="14" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2475" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7948" />
                    <RANKING order="2" place="2" resultid="9497" />
                    <RANKING order="3" place="3" resultid="3823" />
                    <RANKING order="4" place="4" resultid="3832" />
                    <RANKING order="5" place="5" resultid="7665" />
                    <RANKING order="6" place="6" resultid="3309" />
                    <RANKING order="7" place="-1" resultid="10300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2476" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3224" />
                    <RANKING order="2" place="2" resultid="8637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2477" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7370" />
                    <RANKING order="2" place="2" resultid="9845" />
                    <RANKING order="3" place="3" resultid="7935" />
                    <RANKING order="4" place="4" resultid="7079" />
                    <RANKING order="5" place="5" resultid="9851" />
                    <RANKING order="6" place="6" resultid="3846" />
                    <RANKING order="7" place="7" resultid="8845" />
                    <RANKING order="8" place="8" resultid="8548" />
                    <RANKING order="9" place="9" resultid="9870" />
                    <RANKING order="10" place="10" resultid="10320" />
                    <RANKING order="11" place="11" resultid="7005" />
                    <RANKING order="12" place="12" resultid="6444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2478" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7964" />
                    <RANKING order="2" place="2" resultid="6338" />
                    <RANKING order="3" place="3" resultid="6323" />
                    <RANKING order="4" place="4" resultid="3866" />
                    <RANKING order="5" place="5" resultid="7661" />
                    <RANKING order="6" place="6" resultid="7366" />
                    <RANKING order="7" place="7" resultid="7574" />
                    <RANKING order="8" place="8" resultid="8641" />
                    <RANKING order="9" place="9" resultid="6497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2479" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8292" />
                    <RANKING order="2" place="2" resultid="8305" />
                    <RANKING order="3" place="3" resultid="6582" />
                    <RANKING order="4" place="4" resultid="7902" />
                    <RANKING order="5" place="5" resultid="3259" />
                    <RANKING order="6" place="6" resultid="9360" />
                    <RANKING order="7" place="7" resultid="7656" />
                    <RANKING order="8" place="8" resultid="9412" />
                    <RANKING order="9" place="9" resultid="3286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2480" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6671" />
                    <RANKING order="2" place="2" resultid="10105" />
                    <RANKING order="3" place="3" resultid="8623" />
                    <RANKING order="4" place="4" resultid="6640" />
                    <RANKING order="5" place="5" resultid="3238" />
                    <RANKING order="6" place="6" resultid="7568" />
                    <RANKING order="7" place="-1" resultid="6748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2481" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6606" />
                    <RANKING order="2" place="2" resultid="9121" />
                    <RANKING order="3" place="3" resultid="6358" />
                    <RANKING order="4" place="4" resultid="6411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2482" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8940" />
                    <RANKING order="2" place="2" resultid="7351" />
                    <RANKING order="3" place="3" resultid="6665" />
                    <RANKING order="4" place="4" resultid="6484" />
                    <RANKING order="5" place="5" resultid="9353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2483" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7342" />
                    <RANKING order="2" place="2" resultid="3215" />
                    <RANKING order="3" place="3" resultid="3204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2484" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4579" />
                    <RANKING order="2" place="2" resultid="8772" />
                    <RANKING order="3" place="3" resultid="3653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2485" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8769" />
                    <RANKING order="2" place="2" resultid="6625" />
                    <RANKING order="3" place="3" resultid="7980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2486" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2487" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2488" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2489" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2490" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10765" daytime="10:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10766" daytime="10:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10767" daytime="10:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10768" daytime="10:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10769" daytime="10:32" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10770" daytime="10:34" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10771" daytime="10:36" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1332" daytime="11:20" gender="M" number="17" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2523" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10647" />
                    <RANKING order="2" place="2" resultid="7084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2524" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7063" />
                    <RANKING order="2" place="2" resultid="3642" />
                    <RANKING order="3" place="3" resultid="3521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2525" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6802" />
                    <RANKING order="2" place="2" resultid="8835" />
                    <RANKING order="3" place="3" resultid="9103" />
                    <RANKING order="4" place="4" resultid="6894" />
                    <RANKING order="5" place="5" resultid="7628" />
                    <RANKING order="6" place="-1" resultid="10260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2526" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9586" />
                    <RANKING order="2" place="2" resultid="9883" />
                    <RANKING order="3" place="3" resultid="8842" />
                    <RANKING order="4" place="4" resultid="6869" />
                    <RANKING order="5" place="5" resultid="8340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2527" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6636" />
                    <RANKING order="2" place="2" resultid="6401" />
                    <RANKING order="3" place="3" resultid="8451" />
                    <RANKING order="4" place="4" resultid="8022" />
                    <RANKING order="5" place="5" resultid="10279" />
                    <RANKING order="6" place="6" resultid="10273" />
                    <RANKING order="7" place="7" resultid="8241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2528" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6984" />
                    <RANKING order="2" place="2" resultid="8202" />
                    <RANKING order="3" place="3" resultid="8206" />
                    <RANKING order="4" place="4" resultid="8217" />
                    <RANKING order="5" place="5" resultid="6741" />
                    <RANKING order="6" place="6" resultid="7623" />
                    <RANKING order="7" place="-1" resultid="8298" />
                    <RANKING order="8" place="-1" resultid="8647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2529" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6526" />
                    <RANKING order="2" place="2" resultid="9450" />
                    <RANKING order="3" place="3" resultid="6344" />
                    <RANKING order="4" place="4" resultid="8499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2530" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7617" />
                    <RANKING order="2" place="2" resultid="8046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2531" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10573" />
                    <RANKING order="2" place="2" resultid="8984" />
                    <RANKING order="3" place="3" resultid="7924" />
                    <RANKING order="4" place="4" resultid="6307" />
                    <RANKING order="5" place="5" resultid="6791" />
                    <RANKING order="6" place="6" resultid="8898" />
                    <RANKING order="7" place="7" resultid="8887" />
                    <RANKING order="8" place="-1" resultid="4561" />
                    <RANKING order="9" place="-1" resultid="7996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2532" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9033" />
                    <RANKING order="2" place="2" resultid="9838" />
                    <RANKING order="3" place="-1" resultid="6529" />
                    <RANKING order="4" place="-1" resultid="8356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2533" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6617" />
                    <RANKING order="2" place="-1" resultid="8924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2534" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6372" />
                    <RANKING order="2" place="-1" resultid="7974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2535" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2536" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2537" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2538" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10791" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10792" daytime="11:27" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10793" daytime="11:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10794" daytime="11:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10795" daytime="11:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10796" daytime="11:43" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1226" daytime="09:00" gender="F" number="10" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2411" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3822" />
                    <RANKING order="2" place="2" resultid="10299" />
                    <RANKING order="3" place="3" resultid="10555" />
                    <RANKING order="4" place="4" resultid="9496" />
                    <RANKING order="5" place="5" resultid="7947" />
                    <RANKING order="6" place="6" resultid="10125" />
                    <RANKING order="7" place="7" resultid="9439" />
                    <RANKING order="8" place="-1" resultid="7664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2412" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7759" />
                    <RANKING order="2" place="-1" resultid="11061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2413" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6783" />
                    <RANKING order="2" place="2" resultid="9346" />
                    <RANKING order="3" place="-1" resultid="8914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2414" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6322" />
                    <RANKING order="2" place="2" resultid="7963" />
                    <RANKING order="3" place="3" resultid="9092" />
                    <RANKING order="4" place="4" resultid="10087" />
                    <RANKING order="5" place="5" resultid="3865" />
                    <RANKING order="6" place="6" resultid="6878" />
                    <RANKING order="7" place="7" resultid="7660" />
                    <RANKING order="8" place="8" resultid="8266" />
                    <RANKING order="9" place="9" resultid="9391" />
                    <RANKING order="10" place="10" resultid="8850" />
                    <RANKING order="11" place="11" resultid="8026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2415" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8955" />
                    <RANKING order="2" place="2" resultid="6587" />
                    <RANKING order="3" place="3" resultid="7655" />
                    <RANKING order="4" place="4" resultid="3258" />
                    <RANKING order="5" place="5" resultid="9359" />
                    <RANKING order="6" place="-1" resultid="6989" />
                    <RANKING order="7" place="-1" resultid="8304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2416" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7355" />
                    <RANKING order="2" place="2" resultid="8960" />
                    <RANKING order="3" place="3" resultid="10104" />
                    <RANKING order="4" place="4" resultid="6676" />
                    <RANKING order="5" place="5" resultid="6639" />
                    <RANKING order="6" place="6" resultid="3237" />
                    <RANKING order="7" place="7" resultid="7567" />
                    <RANKING order="8" place="8" resultid="3264" />
                    <RANKING order="9" place="-1" resultid="6747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2417" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6605" />
                    <RANKING order="2" place="2" resultid="6289" />
                    <RANKING order="3" place="3" resultid="6357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2418" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8930" />
                    <RANKING order="2" place="2" resultid="8088" />
                    <RANKING order="3" place="3" resultid="6664" />
                    <RANKING order="4" place="4" resultid="9112" />
                    <RANKING order="5" place="5" resultid="6483" />
                    <RANKING order="6" place="6" resultid="8779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2419" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7341" />
                    <RANKING order="2" place="2" resultid="6683" />
                    <RANKING order="3" place="3" resultid="3214" />
                    <RANKING order="4" place="4" resultid="9604" />
                    <RANKING order="5" place="5" resultid="3203" />
                    <RANKING order="6" place="6" resultid="6455" />
                    <RANKING order="7" place="7" resultid="10606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2420" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4578" />
                    <RANKING order="2" place="2" resultid="9069" />
                    <RANKING order="3" place="3" resultid="3652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2421" agemax="74" agemin="70" name="Kat J 70-74" />
                <AGEGROUP agegroupid="2422" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2423" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2424" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2425" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2426" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10734" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10735" daytime="09:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10736" daytime="09:03" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10737" daytime="09:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10738" daytime="09:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10739" daytime="09:07" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1242" daytime="09:09" gender="M" number="11" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2427" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10312" />
                    <RANKING order="2" place="2" resultid="8416" />
                    <RANKING order="3" place="3" resultid="10955" />
                    <RANKING order="4" place="4" resultid="10646" />
                    <RANKING order="5" place="5" resultid="10115" />
                    <RANKING order="6" place="-1" resultid="3624" />
                    <RANKING order="7" place="-1" resultid="7146" />
                    <RANKING order="8" place="-1" resultid="9830" />
                    <RANKING order="9" place="-1" resultid="10306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2428" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7602" />
                    <RANKING order="2" place="2" resultid="6297" />
                    <RANKING order="3" place="3" resultid="9910" />
                    <RANKING order="4" place="-1" resultid="9400" />
                    <RANKING order="5" place="-1" resultid="9417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2429" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6601" />
                    <RANKING order="2" place="2" resultid="6893" />
                    <RANKING order="3" place="3" resultid="6558" />
                    <RANKING order="4" place="4" resultid="9891" />
                    <RANKING order="5" place="5" resultid="3877" />
                    <RANKING order="6" place="6" resultid="6882" />
                    <RANKING order="7" place="7" resultid="7093" />
                    <RANKING order="8" place="8" resultid="8858" />
                    <RANKING order="9" place="9" resultid="6957" />
                    <RANKING order="10" place="10" resultid="9797" />
                    <RANKING order="11" place="11" resultid="10948" />
                    <RANKING order="12" place="12" resultid="3891" />
                    <RANKING order="13" place="13" resultid="6055" />
                    <RANKING order="14" place="14" resultid="9819" />
                    <RANKING order="15" place="-1" resultid="8589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2430" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8652" />
                    <RANKING order="2" place="2" resultid="9882" />
                    <RANKING order="3" place="3" resultid="9629" />
                    <RANKING order="4" place="4" resultid="8442" />
                    <RANKING order="5" place="5" resultid="8976" />
                    <RANKING order="6" place="6" resultid="9435" />
                    <RANKING order="7" place="7" resultid="6520" />
                    <RANKING order="8" place="8" resultid="9428" />
                    <RANKING order="9" place="9" resultid="8339" />
                    <RANKING order="10" place="10" resultid="6509" />
                    <RANKING order="11" place="11" resultid="3273" />
                    <RANKING order="12" place="-1" resultid="3250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2431" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6777" />
                    <RANKING order="2" place="2" resultid="10238" />
                    <RANKING order="3" place="3" resultid="8054" />
                    <RANKING order="4" place="4" resultid="9923" />
                    <RANKING order="5" place="5" resultid="8017" />
                    <RANKING order="6" place="6" resultid="9096" />
                    <RANKING order="7" place="7" resultid="8564" />
                    <RANKING order="8" place="8" resultid="8012" />
                    <RANKING order="9" place="9" resultid="10254" />
                    <RANKING order="10" place="10" resultid="8463" />
                    <RANKING order="11" place="11" resultid="7670" />
                    <RANKING order="12" place="-1" resultid="8489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2432" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3788" />
                    <RANKING order="2" place="2" resultid="8646" />
                    <RANKING order="3" place="3" resultid="8199" />
                    <RANKING order="4" place="4" resultid="7415" />
                    <RANKING order="5" place="5" resultid="10082" />
                    <RANKING order="6" place="6" resultid="8252" />
                    <RANKING order="7" place="7" resultid="4569" />
                    <RANKING order="8" place="8" resultid="3302" />
                    <RANKING order="9" place="9" resultid="8425" />
                    <RANKING order="10" place="10" resultid="9406" />
                    <RANKING order="11" place="11" resultid="3887" />
                    <RANKING order="12" place="-1" resultid="6992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2433" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10163" />
                    <RANKING order="2" place="2" resultid="8520" />
                    <RANKING order="3" place="3" resultid="3657" />
                    <RANKING order="4" place="4" resultid="6525" />
                    <RANKING order="5" place="-1" resultid="6436" />
                    <RANKING order="6" place="-1" resultid="7584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2434" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7746" />
                    <RANKING order="2" place="2" resultid="9917" />
                    <RANKING order="3" place="3" resultid="6690" />
                    <RANKING order="4" place="4" resultid="7634" />
                    <RANKING order="5" place="5" resultid="9106" />
                    <RANKING order="6" place="6" resultid="10617" />
                    <RANKING order="7" place="7" resultid="6761" />
                    <RANKING order="8" place="8" resultid="8776" />
                    <RANKING order="9" place="9" resultid="7391" />
                    <RANKING order="10" place="10" resultid="8512" />
                    <RANKING order="11" place="-1" resultid="9342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2435" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10330" />
                    <RANKING order="2" place="2" resultid="8983" />
                    <RANKING order="3" place="3" resultid="7384" />
                    <RANKING order="4" place="4" resultid="6790" />
                    <RANKING order="5" place="5" resultid="7526" />
                    <RANKING order="6" place="6" resultid="6380" />
                    <RANKING order="7" place="7" resultid="7995" />
                    <RANKING order="8" place="8" resultid="4560" />
                    <RANKING order="9" place="9" resultid="6503" />
                    <RANKING order="10" place="10" resultid="6752" />
                    <RANKING order="11" place="-1" resultid="8628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2436" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8459" />
                    <RANKING order="2" place="2" resultid="8063" />
                    <RANKING order="3" place="3" resultid="9032" />
                    <RANKING order="4" place="4" resultid="8990" />
                    <RANKING order="5" place="5" resultid="8381" />
                    <RANKING order="6" place="6" resultid="9837" />
                    <RANKING order="7" place="7" resultid="8786" />
                    <RANKING order="8" place="8" resultid="9056" />
                    <RANKING order="9" place="9" resultid="3278" />
                    <RANKING order="10" place="10" resultid="8355" />
                    <RANKING order="11" place="-1" resultid="7912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2437" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8794" />
                    <RANKING order="2" place="2" resultid="7375" />
                    <RANKING order="3" place="3" resultid="8579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2438" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9062" />
                    <RANKING order="2" place="2" resultid="8432" />
                    <RANKING order="3" place="3" resultid="7973" />
                    <RANKING order="4" place="4" resultid="8314" />
                    <RANKING order="5" place="-1" resultid="8346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2439" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9077" />
                    <RANKING order="2" place="2" resultid="7750" />
                    <RANKING order="3" place="-1" resultid="8543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2440" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2441" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2442" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10740" daytime="09:09" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10741" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10742" daytime="09:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10743" daytime="09:13" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10744" daytime="09:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10745" daytime="09:16" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10746" daytime="09:17" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10747" daytime="09:18" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10748" daytime="09:19" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10749" daytime="09:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10750" daytime="09:21" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10751" daytime="09:23" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="10:38" gender="M" number="15" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2491" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7083" />
                    <RANKING order="2" place="2" resultid="10313" />
                    <RANKING order="3" place="3" resultid="8417" />
                    <RANKING order="4" place="4" resultid="10956" />
                    <RANKING order="5" place="5" resultid="10263" />
                    <RANKING order="6" place="6" resultid="7597" />
                    <RANKING order="7" place="7" resultid="6475" />
                    <RANKING order="8" place="8" resultid="10231" />
                    <RANKING order="9" place="9" resultid="3851" />
                    <RANKING order="10" place="-1" resultid="7147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2492" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7591" />
                    <RANKING order="2" place="2" resultid="6331" />
                    <RANKING order="3" place="3" resultid="7013" />
                    <RANKING order="4" place="4" resultid="8469" />
                    <RANKING order="5" place="5" resultid="10293" />
                    <RANKING order="6" place="6" resultid="8437" />
                    <RANKING order="7" place="7" resultid="7740" />
                    <RANKING order="8" place="8" resultid="6850" />
                    <RANKING order="9" place="9" resultid="3839" />
                    <RANKING order="10" place="10" resultid="9911" />
                    <RANKING order="11" place="11" resultid="7132" />
                    <RANKING order="12" place="12" resultid="6920" />
                    <RANKING order="13" place="13" resultid="3884" />
                    <RANKING order="14" place="-1" resultid="6861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2493" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6799" />
                    <RANKING order="2" place="2" resultid="9225" />
                    <RANKING order="3" place="3" resultid="8968" />
                    <RANKING order="4" place="4" resultid="3878" />
                    <RANKING order="5" place="5" resultid="8553" />
                    <RANKING order="6" place="6" resultid="9876" />
                    <RANKING order="7" place="7" resultid="7153" />
                    <RANKING order="8" place="8" resultid="9892" />
                    <RANKING order="9" place="9" resultid="6883" />
                    <RANKING order="10" place="10" resultid="8590" />
                    <RANKING order="11" place="11" resultid="8859" />
                    <RANKING order="12" place="12" resultid="9443" />
                    <RANKING order="13" place="13" resultid="3827" />
                    <RANKING order="14" place="14" resultid="9798" />
                    <RANKING order="15" place="15" resultid="10949" />
                    <RANKING order="16" place="16" resultid="6056" />
                    <RANKING order="17" place="17" resultid="10569" />
                    <RANKING order="18" place="-1" resultid="6958" />
                    <RANKING order="19" place="-1" resultid="7612" />
                    <RANKING order="20" place="-1" resultid="8456" />
                    <RANKING order="21" place="-1" resultid="8834" />
                    <RANKING order="22" place="-1" resultid="9898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2494" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6396" />
                    <RANKING order="2" place="2" resultid="8443" />
                    <RANKING order="3" place="3" resultid="8907" />
                    <RANKING order="4" place="4" resultid="6659" />
                    <RANKING order="5" place="5" resultid="8328" />
                    <RANKING order="6" place="6" resultid="3189" />
                    <RANKING order="7" place="7" resultid="9436" />
                    <RANKING order="8" place="8" resultid="6888" />
                    <RANKING order="9" place="9" resultid="8574" />
                    <RANKING order="10" place="10" resultid="6899" />
                    <RANKING order="11" place="11" resultid="7639" />
                    <RANKING order="12" place="12" resultid="9614" />
                    <RANKING order="13" place="13" resultid="8526" />
                    <RANKING order="14" place="14" resultid="8363" />
                    <RANKING order="15" place="15" resultid="7019" />
                    <RANKING order="16" place="16" resultid="6510" />
                    <RANKING order="17" place="17" resultid="6998" />
                    <RANKING order="18" place="18" resultid="8607" />
                    <RANKING order="19" place="19" resultid="10660" />
                    <RANKING order="20" place="20" resultid="3274" />
                    <RANKING order="21" place="-1" resultid="9396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2495" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7645" />
                    <RANKING order="2" place="2" resultid="8078" />
                    <RANKING order="3" place="3" resultid="10239" />
                    <RANKING order="4" place="4" resultid="8259" />
                    <RANKING order="5" place="5" resultid="9382" />
                    <RANKING order="6" place="6" resultid="7157" />
                    <RANKING order="7" place="7" resultid="8248" />
                    <RANKING order="8" place="8" resultid="6577" />
                    <RANKING order="9" place="9" resultid="8018" />
                    <RANKING order="10" place="10" resultid="8565" />
                    <RANKING order="11" place="11" resultid="8594" />
                    <RANKING order="12" place="12" resultid="8240" />
                    <RANKING order="13" place="13" resultid="8618" />
                    <RANKING order="14" place="14" resultid="8013" />
                    <RANKING order="15" place="15" resultid="8490" />
                    <RANKING order="16" place="16" resultid="7827" />
                    <RANKING order="17" place="17" resultid="3856" />
                    <RANKING order="18" place="18" resultid="8464" />
                    <RANKING order="19" place="19" resultid="7671" />
                    <RANKING order="20" place="-1" resultid="6652" />
                    <RANKING order="21" place="-1" resultid="6969" />
                    <RANKING order="22" place="-1" resultid="7795" />
                    <RANKING order="23" place="-1" resultid="8466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2496" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8540" />
                    <RANKING order="2" place="2" resultid="7782" />
                    <RANKING order="3" place="3" resultid="6979" />
                    <RANKING order="4" place="4" resultid="10168" />
                    <RANKING order="5" place="5" resultid="10083" />
                    <RANKING order="6" place="6" resultid="4570" />
                    <RANKING order="7" place="7" resultid="8426" />
                    <RANKING order="8" place="8" resultid="3303" />
                    <RANKING order="9" place="9" resultid="10655" />
                    <RANKING order="10" place="10" resultid="8477" />
                    <RANKING order="11" place="11" resultid="7022" />
                    <RANKING order="12" place="-1" resultid="3295" />
                    <RANKING order="13" place="-1" resultid="7411" />
                    <RANKING order="14" place="-1" resultid="8615" />
                    <RANKING order="15" place="-1" resultid="9814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2497" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8521" />
                    <RANKING order="2" place="2" resultid="6284" />
                    <RANKING order="3" place="3" resultid="6429" />
                    <RANKING order="4" place="4" resultid="10578" />
                    <RANKING order="5" place="5" resultid="8320" />
                    <RANKING order="6" place="6" resultid="7585" />
                    <RANKING order="7" place="7" resultid="8600" />
                    <RANKING order="8" place="8" resultid="6631" />
                    <RANKING order="9" place="9" resultid="7607" />
                    <RANKING order="10" place="10" resultid="7535" />
                    <RANKING order="11" place="11" resultid="10284" />
                    <RANKING order="12" place="12" resultid="9809" />
                    <RANKING order="13" place="-1" resultid="6437" />
                    <RANKING order="14" place="-1" resultid="9449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2498" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8505" />
                    <RANKING order="2" place="2" resultid="9620" />
                    <RANKING order="3" place="3" resultid="9918" />
                    <RANKING order="4" place="4" resultid="7635" />
                    <RANKING order="5" place="5" resultid="8951" />
                    <RANKING order="6" place="6" resultid="6762" />
                    <RANKING order="7" place="7" resultid="6405" />
                    <RANKING order="8" place="8" resultid="8513" />
                    <RANKING order="9" place="9" resultid="6350" />
                    <RANKING order="10" place="-1" resultid="6691" />
                    <RANKING order="11" place="-1" resultid="9117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2499" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8532" />
                    <RANKING order="2" place="2" resultid="9927" />
                    <RANKING order="3" place="3" resultid="7385" />
                    <RANKING order="4" place="4" resultid="10267" />
                    <RANKING order="5" place="5" resultid="6381" />
                    <RANKING order="6" place="6" resultid="6504" />
                    <RANKING order="7" place="7" resultid="8897" />
                    <RANKING order="8" place="8" resultid="7106" />
                    <RANKING order="9" place="9" resultid="6753" />
                    <RANKING order="10" place="-1" resultid="6772" />
                    <RANKING order="11" place="-1" resultid="7527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2500" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8333" />
                    <RANKING order="2" place="2" resultid="8064" />
                    <RANKING order="3" place="3" resultid="8782" />
                    <RANKING order="4" place="4" resultid="7552" />
                    <RANKING order="5" place="5" resultid="9057" />
                    <RANKING order="6" place="6" resultid="3279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2501" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8923" />
                    <RANKING order="2" place="2" resultid="6616" />
                    <RANKING order="3" place="3" resultid="7775" />
                    <RANKING order="4" place="4" resultid="8580" />
                    <RANKING order="5" place="5" resultid="7988" />
                    <RANKING order="6" place="-1" resultid="8795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2502" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8765" />
                    <RANKING order="2" place="2" resultid="6644" />
                    <RANKING order="3" place="3" resultid="8315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2503" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7751" />
                    <RANKING order="2" place="2" resultid="8351" />
                    <RANKING order="3" place="3" resultid="11056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2504" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3245" />
                    <RANKING order="2" place="2" resultid="3161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2505" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2506" agemax="99" agemin="95" name="Kat O 95-99">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="8882" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10772" daytime="10:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10773" daytime="10:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10774" daytime="10:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10775" daytime="10:46" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10776" daytime="10:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10777" daytime="10:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10778" daytime="10:52" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10779" daytime="10:54" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10780" daytime="10:55" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10781" daytime="10:57" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10782" daytime="10:59" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10783" daytime="11:00" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="10784" daytime="11:02" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="10785" daytime="11:03" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="10786" daytime="11:05" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="10787" daytime="11:06" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="10788" daytime="11:08" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2017-06-17" daytime="16:00" endtime="20:43" name="Blok IV" number="4" warmupfrom="14:30" warmupuntil="15:50">
          <EVENTS>
            <EVENT eventid="1422" daytime="16:46" gender="M" number="23" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2587" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10314" />
                    <RANKING order="2" place="2" resultid="7085" />
                    <RANKING order="3" place="3" resultid="8418" />
                    <RANKING order="4" place="4" resultid="6846" />
                    <RANKING order="5" place="5" resultid="6389" />
                    <RANKING order="6" place="6" resultid="10957" />
                    <RANKING order="7" place="7" resultid="7598" />
                    <RANKING order="8" place="8" resultid="6476" />
                    <RANKING order="9" place="9" resultid="10233" />
                    <RANKING order="10" place="-1" resultid="7148" />
                    <RANKING order="11" place="-1" resultid="9831" />
                    <RANKING order="12" place="-1" resultid="10308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2588" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7592" />
                    <RANKING order="2" place="2" resultid="8470" />
                    <RANKING order="3" place="3" resultid="6815" />
                    <RANKING order="4" place="4" resultid="7010" />
                    <RANKING order="5" place="5" resultid="6332" />
                    <RANKING order="6" place="6" resultid="6851" />
                    <RANKING order="7" place="7" resultid="7139" />
                    <RANKING order="8" place="8" resultid="6921" />
                    <RANKING order="9" place="9" resultid="7741" />
                    <RANKING order="10" place="10" resultid="7133" />
                    <RANKING order="11" place="11" resultid="3840" />
                    <RANKING order="12" place="12" resultid="9401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2589" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6797" />
                    <RANKING order="2" place="1" resultid="7909" />
                    <RANKING order="3" place="3" resultid="7011" />
                    <RANKING order="4" place="4" resultid="6559" />
                    <RANKING order="5" place="5" resultid="9807" />
                    <RANKING order="6" place="6" resultid="6884" />
                    <RANKING order="7" place="7" resultid="9893" />
                    <RANKING order="8" place="8" resultid="7792" />
                    <RANKING order="9" place="9" resultid="3879" />
                    <RANKING order="10" place="10" resultid="6906" />
                    <RANKING order="11" place="11" resultid="8860" />
                    <RANKING order="12" place="12" resultid="6959" />
                    <RANKING order="13" place="13" resultid="9444" />
                    <RANKING order="14" place="14" resultid="9821" />
                    <RANKING order="15" place="-1" resultid="7094" />
                    <RANKING order="16" place="-1" resultid="7613" />
                    <RANKING order="17" place="-1" resultid="9226" />
                    <RANKING order="18" place="-1" resultid="9899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2590" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9884" />
                    <RANKING order="2" place="2" resultid="8653" />
                    <RANKING order="3" place="3" resultid="6397" />
                    <RANKING order="4" place="4" resultid="6521" />
                    <RANKING order="5" place="5" resultid="10562" />
                    <RANKING order="6" place="6" resultid="8909" />
                    <RANKING order="7" place="7" resultid="6889" />
                    <RANKING order="8" place="8" resultid="6870" />
                    <RANKING order="9" place="9" resultid="10642" />
                    <RANKING order="10" place="10" resultid="6511" />
                    <RANKING order="11" place="11" resultid="6876" />
                    <RANKING order="12" place="12" resultid="6900" />
                    <RANKING order="13" place="13" resultid="8527" />
                    <RANKING order="14" place="14" resultid="9616" />
                    <RANKING order="15" place="15" resultid="8364" />
                    <RANKING order="16" place="16" resultid="10661" />
                    <RANKING order="17" place="-1" resultid="6660" />
                    <RANKING order="18" place="-1" resultid="9397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2591" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6778" />
                    <RANKING order="2" place="2" resultid="8079" />
                    <RANKING order="3" place="3" resultid="9383" />
                    <RANKING order="4" place="4" resultid="6653" />
                    <RANKING order="5" place="5" resultid="8019" />
                    <RANKING order="6" place="6" resultid="8249" />
                    <RANKING order="7" place="7" resultid="8014" />
                    <RANKING order="8" place="8" resultid="3857" />
                    <RANKING order="9" place="9" resultid="10274" />
                    <RANKING order="10" place="10" resultid="7672" />
                    <RANKING order="11" place="-1" resultid="8492" />
                    <RANKING order="12" place="-1" resultid="10160" />
                    <RANKING order="13" place="-1" resultid="8619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2592" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6985" />
                    <RANKING order="2" place="2" resultid="9051" />
                    <RANKING order="3" place="3" resultid="6980" />
                    <RANKING order="4" place="4" resultid="8203" />
                    <RANKING order="5" place="5" resultid="7783" />
                    <RANKING order="6" place="6" resultid="8648" />
                    <RANKING order="7" place="7" resultid="8207" />
                    <RANKING order="8" place="8" resultid="10169" />
                    <RANKING order="9" place="9" resultid="4571" />
                    <RANKING order="10" place="10" resultid="8218" />
                    <RANKING order="11" place="11" resultid="3304" />
                    <RANKING order="12" place="12" resultid="8427" />
                    <RANKING order="13" place="13" resultid="10656" />
                    <RANKING order="14" place="14" resultid="9815" />
                    <RANKING order="15" place="-1" resultid="7024" />
                    <RANKING order="16" place="-1" resultid="8230" />
                    <RANKING order="17" place="-1" resultid="8255" />
                    <RANKING order="18" place="-1" resultid="8616" />
                    <RANKING order="19" place="-1" resultid="9784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2593" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6438" />
                    <RANKING order="2" place="2" resultid="6285" />
                    <RANKING order="3" place="3" resultid="10164" />
                    <RANKING order="4" place="4" resultid="3658" />
                    <RANKING order="5" place="5" resultid="6430" />
                    <RANKING order="6" place="6" resultid="10579" />
                    <RANKING order="7" place="7" resultid="6807" />
                    <RANKING order="8" place="8" resultid="7586" />
                    <RANKING order="9" place="9" resultid="9451" />
                    <RANKING order="10" place="10" resultid="6633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2594" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8506" />
                    <RANKING order="2" place="2" resultid="6692" />
                    <RANKING order="3" place="3" resultid="9621" />
                    <RANKING order="4" place="4" resultid="7618" />
                    <RANKING order="5" place="5" resultid="8514" />
                    <RANKING order="6" place="6" resultid="7942" />
                    <RANKING order="7" place="7" resultid="6351" />
                    <RANKING order="8" place="-1" resultid="7578" />
                    <RANKING order="9" place="-1" resultid="8047" />
                    <RANKING order="10" place="-1" resultid="9379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2595" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8985" />
                    <RANKING order="2" place="2" resultid="6773" />
                    <RANKING order="3" place="3" resultid="7386" />
                    <RANKING order="4" place="4" resultid="6754" />
                    <RANKING order="5" place="-1" resultid="10268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2596" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8783" />
                    <RANKING order="2" place="2" resultid="8334" />
                    <RANKING order="3" place="3" resultid="9058" />
                    <RANKING order="4" place="4" resultid="8382" />
                    <RANKING order="5" place="5" resultid="9839" />
                    <RANKING order="6" place="6" resultid="8787" />
                    <RANKING order="7" place="-1" resultid="6530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2597" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7777" />
                    <RANKING order="2" place="2" resultid="8925" />
                    <RANKING order="3" place="3" resultid="7376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2598" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6374" />
                    <RANKING order="2" place="2" resultid="8210" />
                    <RANKING order="3" place="3" resultid="7975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2599" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="8545" />
                    <RANKING order="2" place="-1" resultid="11057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2600" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2601" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2602" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10825" daytime="16:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10826" daytime="16:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10827" daytime="16:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10828" daytime="16:51" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10829" daytime="16:52" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10830" daytime="16:54" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10831" daytime="16:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10832" daytime="16:56" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10833" daytime="16:57" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10834" daytime="16:58" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10835" daytime="16:59" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10836" daytime="17:00" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="10837" daytime="17:01" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="10838" daytime="17:02" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1376" daytime="16:00" gender="F" number="20" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2539" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9387" />
                    <RANKING order="2" place="2" resultid="9634" />
                    <RANKING order="3" place="3" resultid="10127" />
                    <RANKING order="4" place="4" resultid="7090" />
                    <RANKING order="5" place="5" resultid="3310" />
                    <RANKING order="6" place="6" resultid="3196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2540" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2541" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8376" />
                    <RANKING order="2" place="2" resultid="10295" />
                    <RANKING order="3" place="3" resultid="9846" />
                    <RANKING order="4" place="4" resultid="8915" />
                    <RANKING order="5" place="5" resultid="8612" />
                    <RANKING order="6" place="6" resultid="6592" />
                    <RANKING order="7" place="7" resultid="8846" />
                    <RANKING order="8" place="8" resultid="9500" />
                    <RANKING order="9" place="9" resultid="9871" />
                    <RANKING order="10" place="10" resultid="8662" />
                    <RANKING order="11" place="11" resultid="3847" />
                    <RANKING order="12" place="12" resultid="8484" />
                    <RANKING order="13" place="13" resultid="9852" />
                    <RANKING order="14" place="14" resultid="3873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2542" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6324" />
                    <RANKING order="2" place="2" resultid="8268" />
                    <RANKING order="3" place="3" resultid="7367" />
                    <RANKING order="4" place="4" resultid="8027" />
                    <RANKING order="5" place="5" resultid="9392" />
                    <RANKING order="6" place="6" resultid="6498" />
                    <RANKING order="7" place="7" resultid="8852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2543" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6317" />
                    <RANKING order="2" place="2" resultid="9534" />
                    <RANKING order="3" place="3" resultid="9488" />
                    <RANKING order="4" place="4" resultid="9413" />
                    <RANKING order="5" place="5" resultid="8293" />
                    <RANKING order="6" place="6" resultid="3287" />
                    <RANKING order="7" place="7" resultid="7834" />
                    <RANKING order="8" place="-1" resultid="6583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2544" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3648" />
                    <RANKING order="2" place="2" resultid="8790" />
                    <RANKING order="3" place="3" resultid="8624" />
                    <RANKING order="4" place="4" resultid="10106" />
                    <RANKING order="5" place="5" resultid="3266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2545" agemax="54" agemin="50" name="Kat F 50-54" />
                <AGEGROUP agegroupid="2546" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8941" />
                    <RANKING order="2" place="2" resultid="9354" />
                    <RANKING order="3" place="3" resultid="6492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2547" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9580" />
                    <RANKING order="2" place="2" resultid="10094" />
                    <RANKING order="3" place="3" resultid="7336" />
                    <RANKING order="4" place="4" resultid="8311" />
                    <RANKING order="5" place="5" resultid="7348" />
                    <RANKING order="6" place="6" resultid="9606" />
                    <RANKING order="7" place="7" resultid="7563" />
                    <RANKING order="8" place="8" resultid="10608" />
                    <RANKING order="9" place="-1" resultid="6457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2548" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2549" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8761" />
                    <RANKING order="2" place="2" resultid="6626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2550" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2551" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2552" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2553" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2554" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10803" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10804" daytime="16:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10805" daytime="16:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10806" daytime="16:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10807" daytime="16:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10808" daytime="16:12" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1497" daytime="18:31" gender="F" number="28" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1512" agemax="119" agemin="100" name="Kat A 100-119" />
                <AGEGROUP agegroupid="1513" agemax="159" agemin="120" name="Kat B 120-159">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9904" />
                    <RANKING order="2" place="2" resultid="8675" />
                    <RANKING order="3" place="3" resultid="8676" />
                    <RANKING order="4" place="4" resultid="8867" />
                    <RANKING order="5" place="-1" resultid="9464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1514" agemax="199" agemin="160" name="Kat C 160-199">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1515" agemax="239" agemin="200" name="Kat D 200-239">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6702" />
                    <RANKING order="2" place="2" resultid="9000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1516" agemax="279" agemin="240" name="Kat E 240-279">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8802" />
                    <RANKING order="2" place="2" resultid="7432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="-1" agemin="280" name="Kat F 280 +" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10867" daytime="18:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10868" daytime="18:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1392" daytime="16:15" gender="M" number="21" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2555" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6388" />
                    <RANKING order="2" place="2" resultid="9520" />
                    <RANKING order="3" place="3" resultid="10117" />
                    <RANKING order="4" place="4" resultid="10232" />
                    <RANKING order="5" place="-1" resultid="3626" />
                    <RANKING order="6" place="-1" resultid="10307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2556" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9531" />
                    <RANKING order="2" place="2" resultid="7071" />
                    <RANKING order="3" place="3" resultid="3522" />
                    <RANKING order="4" place="4" resultid="6299" />
                    <RANKING order="5" place="5" resultid="7138" />
                    <RANKING order="6" place="-1" resultid="6857" />
                    <RANKING order="7" place="-1" resultid="8222" />
                    <RANKING order="8" place="-1" resultid="10566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2557" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8370" />
                    <RANKING order="2" place="2" resultid="8604" />
                    <RANKING order="3" place="3" resultid="8969" />
                    <RANKING order="4" place="4" resultid="9877" />
                    <RANKING order="5" place="5" resultid="7791" />
                    <RANKING order="6" place="6" resultid="6905" />
                    <RANKING order="7" place="7" resultid="10612" />
                    <RANKING order="8" place="8" resultid="6303" />
                    <RANKING order="9" place="9" resultid="9799" />
                    <RANKING order="10" place="10" resultid="3828" />
                    <RANKING order="11" place="11" resultid="9820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2558" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8561" />
                    <RANKING order="2" place="2" resultid="8908" />
                    <RANKING order="3" place="3" resultid="9615" />
                    <RANKING order="4" place="4" resultid="6875" />
                    <RANKING order="5" place="5" resultid="6914" />
                    <RANKING order="6" place="6" resultid="3275" />
                    <RANKING order="7" place="7" resultid="3252" />
                    <RANKING order="8" place="-1" resultid="10290" />
                    <RANKING order="9" place="-1" resultid="10561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2559" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8008" />
                    <RANKING order="2" place="2" resultid="8260" />
                    <RANKING order="3" place="3" resultid="6611" />
                    <RANKING order="4" place="4" resultid="8566" />
                    <RANKING order="5" place="5" resultid="10621" />
                    <RANKING order="6" place="6" resultid="8056" />
                    <RANKING order="7" place="7" resultid="8595" />
                    <RANKING order="8" place="8" resultid="10256" />
                    <RANKING order="9" place="9" resultid="6578" />
                    <RANKING order="10" place="10" resultid="8491" />
                    <RANKING order="11" place="11" resultid="3183" />
                    <RANKING order="12" place="12" resultid="9792" />
                    <RANKING order="13" place="-1" resultid="6970" />
                    <RANKING order="14" place="-1" resultid="7796" />
                    <RANKING order="15" place="-1" resultid="10159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2560" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6422" />
                    <RANKING order="2" place="2" resultid="8234" />
                    <RANKING order="3" place="3" resultid="8229" />
                    <RANKING order="4" place="4" resultid="3296" />
                    <RANKING order="5" place="5" resultid="7788" />
                    <RANKING order="6" place="6" resultid="6742" />
                    <RANKING order="7" place="7" resultid="8254" />
                    <RANKING order="8" place="8" resultid="8478" />
                    <RANKING order="9" place="9" resultid="9407" />
                    <RANKING order="10" place="-1" resultid="7023" />
                    <RANKING order="11" place="-1" resultid="6974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2561" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7405" />
                    <RANKING order="2" place="2" resultid="7398" />
                    <RANKING order="3" place="3" resultid="8601" />
                    <RANKING order="4" place="4" resultid="6632" />
                    <RANKING order="5" place="5" resultid="8500" />
                    <RANKING order="6" place="6" resultid="9788" />
                    <RANKING order="7" place="7" resultid="7536" />
                    <RANKING order="8" place="8" resultid="6329" />
                    <RANKING order="9" place="9" resultid="10285" />
                    <RANKING order="10" place="10" resultid="9810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2562" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6537" />
                    <RANKING order="2" place="2" resultid="9626" />
                    <RANKING order="3" place="3" resultid="9108" />
                    <RANKING order="4" place="4" resultid="8920" />
                    <RANKING order="5" place="5" resultid="8952" />
                    <RANKING order="6" place="6" resultid="7392" />
                    <RANKING order="7" place="-1" resultid="7547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2563" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10574" />
                    <RANKING order="2" place="2" resultid="10331" />
                    <RANKING order="3" place="3" resultid="7925" />
                    <RANKING order="4" place="4" resultid="9074" />
                    <RANKING order="5" place="5" resultid="6308" />
                    <RANKING order="6" place="6" resultid="8558" />
                    <RANKING order="7" place="7" resultid="9126" />
                    <RANKING order="8" place="8" resultid="6554" />
                    <RANKING order="9" place="-1" resultid="6382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2564" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8633" />
                    <RANKING order="2" place="2" resultid="8892" />
                    <RANKING order="3" place="3" resultid="8947" />
                    <RANKING order="4" place="4" resultid="7380" />
                    <RANKING order="5" place="5" resultid="8991" />
                    <RANKING order="6" place="6" resultid="3231" />
                    <RANKING order="7" place="-1" resultid="7557" />
                    <RANKING order="8" place="-1" resultid="7913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2565" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7479" />
                    <RANKING order="2" place="2" resultid="7831" />
                    <RANKING order="3" place="3" resultid="7776" />
                    <RANKING order="4" place="4" resultid="7989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2566" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8758" />
                    <RANKING order="2" place="2" resultid="6373" />
                    <RANKING order="3" place="3" resultid="8433" />
                    <RANKING order="4" place="4" resultid="9064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2567" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9078" />
                    <RANKING order="2" place="-1" resultid="8352" />
                    <RANKING order="3" place="-1" resultid="8544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2568" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3246" />
                    <RANKING order="2" place="2" resultid="3162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2569" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2570" agemax="99" agemin="95" name="Kat O 95-99">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7324" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10809" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10810" daytime="16:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10811" daytime="16:21" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10812" daytime="16:23" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10813" daytime="16:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10814" daytime="16:27" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10815" daytime="16:29" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10816" daytime="16:31" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10817" daytime="16:33" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10818" daytime="16:35" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10819" daytime="16:37" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1407" daytime="16:39" gender="F" number="22" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2571" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9490" />
                    <RANKING order="2" place="2" resultid="7949" />
                    <RANKING order="3" place="3" resultid="9635" />
                    <RANKING order="4" place="4" resultid="7679" />
                    <RANKING order="5" place="5" resultid="3833" />
                    <RANKING order="6" place="6" resultid="7666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2572" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2573" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7371" />
                    <RANKING order="2" place="2" resultid="7936" />
                    <RANKING order="3" place="3" resultid="8916" />
                    <RANKING order="4" place="4" resultid="8549" />
                    <RANKING order="5" place="5" resultid="9501" />
                    <RANKING order="6" place="6" resultid="8663" />
                    <RANKING order="7" place="7" resultid="7006" />
                    <RANKING order="8" place="-1" resultid="6784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2574" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7965" />
                    <RANKING order="2" place="2" resultid="6879" />
                    <RANKING order="3" place="3" resultid="9093" />
                    <RANKING order="4" place="4" resultid="6339" />
                    <RANKING order="5" place="5" resultid="10088" />
                    <RANKING order="6" place="6" resultid="9424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2575" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6318" />
                    <RANKING order="2" place="2" resultid="7903" />
                    <RANKING order="3" place="3" resultid="8306" />
                    <RANKING order="4" place="4" resultid="6656" />
                    <RANKING order="5" place="-1" resultid="6990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2576" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7357" />
                    <RANKING order="2" place="2" resultid="6672" />
                    <RANKING order="3" place="3" resultid="8962" />
                    <RANKING order="4" place="4" resultid="6677" />
                    <RANKING order="5" place="5" resultid="10107" />
                    <RANKING order="6" place="6" resultid="6641" />
                    <RANKING order="7" place="-1" resultid="6749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2577" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6607" />
                    <RANKING order="2" place="2" resultid="8072" />
                    <RANKING order="3" place="3" resultid="6412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2578" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8932" />
                    <RANKING order="2" place="2" resultid="6666" />
                    <RANKING order="3" place="3" resultid="9355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2579" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7343" />
                    <RANKING order="2" place="2" resultid="10095" />
                    <RANKING order="3" place="3" resultid="6685" />
                    <RANKING order="4" place="4" resultid="8312" />
                    <RANKING order="5" place="5" resultid="3205" />
                    <RANKING order="6" place="-1" resultid="3216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2580" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4580" />
                    <RANKING order="2" place="2" resultid="3654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2581" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2582" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2583" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2584" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2585" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2586" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10820" daytime="16:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10821" daytime="16:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10822" daytime="16:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10823" daytime="16:43" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10824" daytime="16:45" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1437" daytime="17:03" gender="F" number="24" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2603" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3824" />
                    <RANKING order="2" place="2" resultid="10556" />
                    <RANKING order="3" place="3" resultid="3834" />
                    <RANKING order="4" place="-1" resultid="10128" />
                    <RANKING order="5" place="-1" resultid="10301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2604" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2605" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6785" />
                    <RANKING order="2" place="2" resultid="9347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2606" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3867" />
                    <RANKING order="2" place="2" resultid="7966" />
                    <RANKING order="3" place="3" resultid="10089" />
                    <RANKING order="4" place="4" resultid="9094" />
                    <RANKING order="5" place="5" resultid="8853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2607" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8956" />
                    <RANKING order="2" place="2" resultid="7159" />
                    <RANKING order="3" place="3" resultid="8829" />
                    <RANKING order="4" place="4" resultid="6588" />
                    <RANKING order="5" place="5" resultid="7657" />
                    <RANKING order="6" place="6" resultid="3260" />
                    <RANKING order="7" place="7" resultid="9361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2608" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8963" />
                    <RANKING order="2" place="2" resultid="6678" />
                    <RANKING order="3" place="3" resultid="7569" />
                    <RANKING order="4" place="4" resultid="3267" />
                    <RANKING order="5" place="-1" resultid="6750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2609" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6608" />
                    <RANKING order="2" place="2" resultid="6291" />
                    <RANKING order="3" place="3" resultid="6359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2610" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8089" />
                    <RANKING order="2" place="2" resultid="9113" />
                    <RANKING order="3" place="3" resultid="8933" />
                    <RANKING order="4" place="4" resultid="6485" />
                    <RANKING order="5" place="5" resultid="9597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2611" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3217" />
                    <RANKING order="2" place="2" resultid="6458" />
                    <RANKING order="3" place="-1" resultid="7337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2612" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2613" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2614" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2615" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2616" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2617" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2618" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10839" daytime="17:03" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10840" daytime="17:07" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10841" daytime="17:09" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10842" daytime="17:11" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1467" daytime="17:31" gender="F" number="26" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2635" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6391" />
                    <RANKING order="2" place="2" resultid="9491" />
                    <RANKING order="3" place="3" resultid="7667" />
                    <RANKING order="4" place="4" resultid="3311" />
                    <RANKING order="5" place="-1" resultid="7950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2636" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3225" />
                    <RANKING order="2" place="2" resultid="3512" />
                    <RANKING order="3" place="-1" resultid="3634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2637" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7372" />
                    <RANKING order="2" place="2" resultid="7080" />
                    <RANKING order="3" place="3" resultid="7937" />
                    <RANKING order="4" place="4" resultid="9861" />
                    <RANKING order="5" place="5" resultid="8550" />
                    <RANKING order="6" place="6" resultid="9853" />
                    <RANKING order="7" place="7" resultid="9872" />
                    <RANKING order="8" place="8" resultid="6445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2638" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6340" />
                    <RANKING order="2" place="2" resultid="3868" />
                    <RANKING order="3" place="3" resultid="8642" />
                    <RANKING order="4" place="4" resultid="6499" />
                    <RANKING order="5" place="5" resultid="9425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2639" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7904" />
                    <RANKING order="2" place="2" resultid="6584" />
                    <RANKING order="3" place="3" resultid="8294" />
                    <RANKING order="4" place="4" resultid="8307" />
                    <RANKING order="5" place="5" resultid="3261" />
                    <RANKING order="6" place="6" resultid="9362" />
                    <RANKING order="7" place="7" resultid="6767" />
                    <RANKING order="8" place="8" resultid="6657" />
                    <RANKING order="9" place="-1" resultid="3288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2640" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8625" />
                    <RANKING order="2" place="2" resultid="3239" />
                    <RANKING order="3" place="3" resultid="7570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2641" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9122" />
                    <RANKING order="2" place="2" resultid="6360" />
                    <RANKING order="3" place="3" resultid="6413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2642" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7352" />
                    <RANKING order="2" place="2" resultid="8942" />
                    <RANKING order="3" place="3" resultid="6667" />
                    <RANKING order="4" place="4" resultid="6486" />
                    <RANKING order="5" place="5" resultid="6450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2643" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7344" />
                    <RANKING order="2" place="2" resultid="3206" />
                    <RANKING order="3" place="3" resultid="9607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2644" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4581" />
                    <RANKING order="2" place="2" resultid="8773" />
                    <RANKING order="3" place="3" resultid="8571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2645" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2646" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2647" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2648" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2649" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2650" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10851" daytime="17:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10852" daytime="17:37" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10853" daytime="17:41" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10854" daytime="17:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10855" daytime="17:48" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1452" daytime="17:13" gender="M" number="25" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2619" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10648" />
                    <RANKING order="2" place="2" resultid="8419" />
                    <RANKING order="3" place="3" resultid="10958" />
                    <RANKING order="4" place="-1" resultid="3627" />
                    <RANKING order="5" place="-1" resultid="9832" />
                    <RANKING order="6" place="-1" resultid="10118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2620" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7603" />
                    <RANKING order="2" place="2" resultid="6300" />
                    <RANKING order="3" place="3" resultid="9912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2621" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6602" />
                    <RANKING order="2" place="2" resultid="6895" />
                    <RANKING order="3" place="3" resultid="6560" />
                    <RANKING order="4" place="4" resultid="9894" />
                    <RANKING order="5" place="5" resultid="9800" />
                    <RANKING order="6" place="6" resultid="10950" />
                    <RANKING order="7" place="7" resultid="8861" />
                    <RANKING order="8" place="8" resultid="3892" />
                    <RANKING order="9" place="9" resultid="6057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2622" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9885" />
                    <RANKING order="2" place="2" resultid="8654" />
                    <RANKING order="3" place="3" resultid="9630" />
                    <RANKING order="4" place="4" resultid="8444" />
                    <RANKING order="5" place="5" resultid="8977" />
                    <RANKING order="6" place="6" resultid="9429" />
                    <RANKING order="7" place="7" resultid="8341" />
                    <RANKING order="8" place="8" resultid="6512" />
                    <RANKING order="9" place="9" resultid="3253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2623" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6779" />
                    <RANKING order="2" place="2" resultid="10240" />
                    <RANKING order="3" place="3" resultid="9515" />
                    <RANKING order="4" place="4" resultid="9924" />
                    <RANKING order="5" place="5" resultid="8057" />
                    <RANKING order="6" place="6" resultid="9098" />
                    <RANKING order="7" place="7" resultid="8023" />
                    <RANKING order="8" place="8" resultid="6572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2624" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3789" />
                    <RANKING order="2" place="2" resultid="8200" />
                    <RANKING order="3" place="3" resultid="7416" />
                    <RANKING order="4" place="4" resultid="9408" />
                    <RANKING order="5" place="-1" resultid="6993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2625" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10165" />
                    <RANKING order="2" place="2" resultid="8522" />
                    <RANKING order="3" place="3" resultid="10580" />
                    <RANKING order="4" place="4" resultid="7406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2626" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7747" />
                    <RANKING order="2" place="2" resultid="9919" />
                    <RANKING order="3" place="3" resultid="6693" />
                    <RANKING order="4" place="4" resultid="7636" />
                    <RANKING order="5" place="5" resultid="9109" />
                    <RANKING order="6" place="6" resultid="6763" />
                    <RANKING order="7" place="7" resultid="10618" />
                    <RANKING order="8" place="8" resultid="8777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2627" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8533" />
                    <RANKING order="2" place="2" resultid="4562" />
                    <RANKING order="3" place="3" resultid="6792" />
                    <RANKING order="4" place="4" resultid="7997" />
                    <RANKING order="5" place="5" resultid="6505" />
                    <RANKING order="6" place="6" resultid="7528" />
                    <RANKING order="7" place="7" resultid="8629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2628" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8460" />
                    <RANKING order="2" place="2" resultid="8065" />
                    <RANKING order="3" place="3" resultid="9034" />
                    <RANKING order="4" place="4" resultid="8383" />
                    <RANKING order="5" place="5" resultid="8992" />
                    <RANKING order="6" place="6" resultid="3280" />
                    <RANKING order="7" place="-1" resultid="6531" />
                    <RANKING order="8" place="-1" resultid="7914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2629" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8796" />
                    <RANKING order="2" place="2" resultid="8581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2630" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9065" />
                    <RANKING order="2" place="2" resultid="8434" />
                    <RANKING order="3" place="3" resultid="8347" />
                    <RANKING order="4" place="4" resultid="8316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2631" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9079" />
                    <RANKING order="2" place="2" resultid="7752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2632" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2633" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2634" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10843" daytime="17:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10844" daytime="17:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10845" daytime="17:19" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10846" daytime="17:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10847" daytime="17:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10848" daytime="17:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10849" daytime="17:27" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10850" daytime="17:29" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1482" daytime="17:52" gender="M" number="27" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2651" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7086" />
                    <RANKING order="2" place="2" resultid="6477" />
                    <RANKING order="3" place="3" resultid="7599" />
                    <RANKING order="4" place="-1" resultid="10264" />
                    <RANKING order="5" place="-1" resultid="10315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2652" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7593" />
                    <RANKING order="2" place="2" resultid="3643" />
                    <RANKING order="3" place="3" resultid="8438" />
                    <RANKING order="4" place="4" resultid="7064" />
                    <RANKING order="5" place="5" resultid="6852" />
                    <RANKING order="6" place="6" resultid="7742" />
                    <RANKING order="7" place="7" resultid="6862" />
                    <RANKING order="8" place="8" resultid="3841" />
                    <RANKING order="9" place="9" resultid="9913" />
                    <RANKING order="10" place="10" resultid="7134" />
                    <RANKING order="11" place="-1" resultid="7014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2653" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8554" />
                    <RANKING order="2" place="2" resultid="7154" />
                    <RANKING order="3" place="3" resultid="8836" />
                    <RANKING order="4" place="4" resultid="8371" />
                    <RANKING order="5" place="5" resultid="8591" />
                    <RANKING order="6" place="6" resultid="6960" />
                    <RANKING order="7" place="7" resultid="7614" />
                    <RANKING order="8" place="8" resultid="10951" />
                    <RANKING order="9" place="9" resultid="6058" />
                    <RANKING order="10" place="-1" resultid="8457" />
                    <RANKING order="11" place="-1" resultid="8970" />
                    <RANKING order="12" place="-1" resultid="10570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2654" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9587" />
                    <RANKING order="2" place="2" resultid="6398" />
                    <RANKING order="3" place="3" resultid="8445" />
                    <RANKING order="4" place="4" resultid="8575" />
                    <RANKING order="5" place="5" resultid="6890" />
                    <RANKING order="6" place="6" resultid="8329" />
                    <RANKING order="7" place="7" resultid="7640" />
                    <RANKING order="8" place="8" resultid="6871" />
                    <RANKING order="9" place="9" resultid="8528" />
                    <RANKING order="10" place="10" resultid="8342" />
                    <RANKING order="11" place="11" resultid="8365" />
                    <RANKING order="12" place="12" resultid="8608" />
                    <RANKING order="13" place="13" resultid="10662" />
                    <RANKING order="14" place="-1" resultid="3276" />
                    <RANKING order="15" place="-1" resultid="9631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2655" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8080" />
                    <RANKING order="2" place="2" resultid="7646" />
                    <RANKING order="3" place="3" resultid="8261" />
                    <RANKING order="4" place="4" resultid="9384" />
                    <RANKING order="5" place="5" resultid="6579" />
                    <RANKING order="6" place="6" resultid="8242" />
                    <RANKING order="7" place="7" resultid="8567" />
                    <RANKING order="8" place="8" resultid="10257" />
                    <RANKING order="9" place="9" resultid="7828" />
                    <RANKING order="10" place="10" resultid="3858" />
                    <RANKING order="11" place="11" resultid="7673" />
                    <RANKING order="12" place="12" resultid="10622" />
                    <RANKING order="13" place="-1" resultid="7797" />
                    <RANKING order="14" place="-1" resultid="8009" />
                    <RANKING order="15" place="-1" resultid="8467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2656" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8541" />
                    <RANKING order="2" place="2" resultid="7784" />
                    <RANKING order="3" place="3" resultid="8649" />
                    <RANKING order="4" place="4" resultid="7412" />
                    <RANKING order="5" place="5" resultid="8299" />
                    <RANKING order="6" place="6" resultid="4572" />
                    <RANKING order="7" place="7" resultid="8428" />
                    <RANKING order="8" place="8" resultid="3305" />
                    <RANKING order="9" place="9" resultid="8479" />
                    <RANKING order="10" place="-1" resultid="3297" />
                    <RANKING order="11" place="-1" resultid="9816" />
                    <RANKING order="12" place="-1" resultid="10084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2657" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6431" />
                    <RANKING order="2" place="2" resultid="8523" />
                    <RANKING order="3" place="3" resultid="8321" />
                    <RANKING order="4" place="4" resultid="7587" />
                    <RANKING order="5" place="5" resultid="8537" />
                    <RANKING order="6" place="6" resultid="7608" />
                    <RANKING order="7" place="7" resultid="7537" />
                    <RANKING order="8" place="8" resultid="10286" />
                    <RANKING order="9" place="-1" resultid="9452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2658" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8507" />
                    <RANKING order="2" place="2" resultid="9118" />
                    <RANKING order="3" place="3" resultid="6406" />
                    <RANKING order="4" place="4" resultid="8515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2659" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8534" />
                    <RANKING order="2" place="2" resultid="7387" />
                    <RANKING order="3" place="3" resultid="9928" />
                    <RANKING order="4" place="4" resultid="10269" />
                    <RANKING order="5" place="5" resultid="6506" />
                    <RANKING order="6" place="6" resultid="8095" />
                    <RANKING order="7" place="7" resultid="8899" />
                    <RANKING order="8" place="-1" resultid="6383" />
                    <RANKING order="9" place="-1" resultid="7529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2660" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8335" />
                    <RANKING order="2" place="2" resultid="7553" />
                    <RANKING order="3" place="3" resultid="8357" />
                    <RANKING order="4" place="4" resultid="3281" />
                    <RANKING order="5" place="5" resultid="3232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2661" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6618" />
                    <RANKING order="2" place="2" resultid="8582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2662" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8766" />
                    <RANKING order="2" place="2" resultid="6645" />
                    <RANKING order="3" place="3" resultid="8348" />
                    <RANKING order="4" place="4" resultid="8317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2663" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7753" />
                    <RANKING order="2" place="-1" resultid="11058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2664" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3247" />
                    <RANKING order="2" place="2" resultid="3163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2665" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2666" agemax="99" agemin="95" name="Kat O 95-99">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8883" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10856" daytime="17:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10857" daytime="17:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10858" daytime="18:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10859" daytime="18:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10860" daytime="18:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10861" daytime="18:13" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10862" daytime="18:16" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10863" daytime="18:19" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10864" daytime="18:22" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10865" daytime="18:25" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10866" daytime="18:27" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1518" daytime="18:37" gender="M" number="29" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1519" agemax="119" agemin="100" name="Kat A 100-119">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1520" agemax="159" agemin="120" name="Kat B 120-159">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6819" />
                    <RANKING order="2" place="2" resultid="7682" />
                    <RANKING order="3" place="3" resultid="6925" />
                    <RANKING order="4" place="4" resultid="8673" />
                    <RANKING order="5" place="5" resultid="3898" />
                    <RANKING order="6" place="6" resultid="9461" />
                    <RANKING order="7" place="7" resultid="6926" />
                    <RANKING order="8" place="-1" resultid="9901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1521" agemax="199" agemin="160" name="Kat C 160-199">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8672" />
                    <RANKING order="2" place="2" resultid="8996" />
                    <RANKING order="3" place="3" resultid="8030" />
                    <RANKING order="4" place="4" resultid="8274" />
                    <RANKING order="5" place="5" resultid="9643" />
                    <RANKING order="6" place="6" resultid="8674" />
                    <RANKING order="7" place="7" resultid="7031" />
                    <RANKING order="8" place="8" resultid="9463" />
                    <RANKING order="9" place="-1" resultid="6820" />
                    <RANKING order="10" place="-1" resultid="7687" />
                    <RANKING order="11" place="-1" resultid="7799" />
                    <RANKING order="12" place="-1" resultid="8387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1522" agemax="239" agemin="200" name="Kat D 200-239">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7436" />
                    <RANKING order="2" place="2" resultid="7686" />
                    <RANKING order="3" place="3" resultid="6703" />
                    <RANKING order="4" place="4" resultid="9131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1523" agemax="279" agemin="240" name="Kat E 240-279">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8998" />
                    <RANKING order="2" place="2" resultid="7433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1524" agemax="-1" agemin="280" name="Kat F 280 +">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8803" />
                    <RANKING order="2" place="2" resultid="9082" />
                    <RANKING order="3" place="3" resultid="8385" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10869" daytime="18:37" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10870" daytime="18:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10871" daytime="18:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10872" daytime="18:48" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1546" daytime="19:16" gender="M" number="31" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2683" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9521" />
                    <RANKING order="2" place="2" resultid="10649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2684" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7604" />
                    <RANKING order="2" place="2" resultid="7065" />
                    <RANKING order="3" place="3" resultid="7072" />
                    <RANKING order="4" place="4" resultid="3523" />
                    <RANKING order="5" place="-1" resultid="6863" />
                    <RANKING order="6" place="-1" resultid="8471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2685" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6803" />
                    <RANKING order="2" place="2" resultid="8837" />
                    <RANKING order="3" place="3" resultid="9104" />
                    <RANKING order="4" place="4" resultid="6896" />
                    <RANKING order="5" place="5" resultid="7630" />
                    <RANKING order="6" place="-1" resultid="3880" />
                    <RANKING order="7" place="-1" resultid="6961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2686" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9588" />
                    <RANKING order="2" place="2" resultid="8843" />
                    <RANKING order="3" place="3" resultid="9430" />
                    <RANKING order="4" place="4" resultid="6916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2687" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7647" />
                    <RANKING order="2" place="2" resultid="8452" />
                    <RANKING order="3" place="3" resultid="9925" />
                    <RANKING order="4" place="4" resultid="6402" />
                    <RANKING order="5" place="5" resultid="6573" />
                    <RANKING order="6" place="6" resultid="8243" />
                    <RANKING order="7" place="7" resultid="8024" />
                    <RANKING order="8" place="8" resultid="10275" />
                    <RANKING order="9" place="-1" resultid="10280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2688" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8235" />
                    <RANKING order="2" place="2" resultid="6743" />
                    <RANKING order="3" place="3" resultid="8300" />
                    <RANKING order="4" place="4" resultid="7624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2689" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6439" />
                    <RANKING order="2" place="2" resultid="6286" />
                    <RANKING order="3" place="3" resultid="7399" />
                    <RANKING order="4" place="4" resultid="6345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2690" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6407" />
                    <RANKING order="2" place="-1" resultid="7579" />
                    <RANKING order="3" place="-1" resultid="7619" />
                    <RANKING order="4" place="-1" resultid="8048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2691" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8986" />
                    <RANKING order="2" place="2" resultid="7926" />
                    <RANKING order="3" place="3" resultid="4563" />
                    <RANKING order="4" place="4" resultid="6309" />
                    <RANKING order="5" place="5" resultid="6793" />
                    <RANKING order="6" place="6" resultid="8900" />
                    <RANKING order="7" place="7" resultid="8888" />
                    <RANKING order="8" place="-1" resultid="7998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2692" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8634" />
                    <RANKING order="2" place="2" resultid="8066" />
                    <RANKING order="3" place="3" resultid="9035" />
                    <RANKING order="4" place="4" resultid="9840" />
                    <RANKING order="5" place="5" resultid="8358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2693" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8926" />
                    <RANKING order="2" place="2" resultid="6619" />
                    <RANKING order="3" place="3" resultid="7990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2694" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2695" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2696" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2697" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2698" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10876" daytime="19:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10877" daytime="19:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10878" daytime="19:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10879" daytime="19:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10880" daytime="19:52" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10881" daytime="19:58" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1525" daytime="18:51" gender="F" number="30" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2667" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7680" />
                    <RANKING order="2" place="2" resultid="3197" />
                    <RANKING order="3" place="-1" resultid="6392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2668" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3226" />
                    <RANKING order="2" place="2" resultid="7761" />
                    <RANKING order="3" place="3" resultid="3513" />
                    <RANKING order="4" place="-1" resultid="3635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2669" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8377" />
                    <RANKING order="2" place="2" resultid="9862" />
                    <RANKING order="3" place="3" resultid="6593" />
                    <RANKING order="4" place="-1" resultid="9348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2670" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6325" />
                    <RANKING order="2" place="2" resultid="8269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2671" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2672" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7358" />
                    <RANKING order="2" place="2" resultid="8791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2673" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6649" />
                    <RANKING order="2" place="2" resultid="6292" />
                    <RANKING order="3" place="-1" resultid="8073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2674" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8090" />
                    <RANKING order="2" place="2" resultid="9598" />
                    <RANKING order="3" place="3" resultid="6493" />
                    <RANKING order="4" place="-1" resultid="6451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2675" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2676" agemax="69" agemin="65" name="Kat I 65-69" />
                <AGEGROUP agegroupid="2677" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2678" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2679" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2680" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2681" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2682" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10873" daytime="18:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10874" daytime="19:01" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10875" daytime="19:09" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2017-06-18" daytime="09:00" name="V Blok" number="5" warmupfrom="07:30" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="1562" daytime="09:00" gender="F" number="32" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2699" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9636" />
                    <RANKING order="2" place="2" resultid="3835" />
                    <RANKING order="3" place="-1" resultid="9639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2700" agemax="29" agemin="25" name="Kat A - 25-29" />
                <AGEGROUP agegroupid="2701" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9502" />
                    <RANKING order="2" place="2" resultid="7007" />
                    <RANKING order="3" place="-1" resultid="6786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2702" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7967" />
                    <RANKING order="2" place="2" resultid="6326" />
                    <RANKING order="3" place="3" resultid="3869" />
                    <RANKING order="4" place="4" resultid="8270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2703" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2704" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8964" />
                    <RANKING order="2" place="2" resultid="6673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2705" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6650" />
                    <RANKING order="2" place="2" resultid="8074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2706" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8934" />
                    <RANKING order="2" place="2" resultid="6452" />
                    <RANKING order="3" place="3" resultid="9599" />
                    <RANKING order="4" place="4" resultid="6494" />
                    <RANKING order="5" place="-1" resultid="6668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2707" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6687" />
                    <RANKING order="2" place="2" resultid="3218" />
                    <RANKING order="3" place="3" resultid="3207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2708" agemax="69" agemin="65" name="Kat I 65-69" />
                <AGEGROUP agegroupid="2709" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8763" />
                    <RANKING order="2" place="2" resultid="6628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2710" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2711" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2712" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2713" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2714" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10882" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10883" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10884" daytime="09:06" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1653" daytime="10:50" number="38" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1668" agemax="119" agemin="100" name="Kat A 100-119">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7032" />
                    <RANKING order="2" place="2" resultid="8677" />
                    <RANKING order="3" place="3" resultid="7097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1669" agemax="159" agemin="120" name="Kat B 120-159">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9908" />
                    <RANKING order="2" place="2" resultid="7688" />
                    <RANKING order="3" place="3" resultid="8865" />
                    <RANKING order="4" place="4" resultid="3895" />
                    <RANKING order="5" place="5" resultid="6595" />
                    <RANKING order="6" place="6" resultid="8678" />
                    <RANKING order="7" place="7" resultid="3317" />
                    <RANKING order="8" place="-1" resultid="9902" />
                    <RANKING order="9" place="-1" resultid="9906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1670" agemax="199" agemin="160" name="Kat C 160-199">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9001" />
                    <RANKING order="2" place="2" resultid="6697" />
                    <RANKING order="3" place="3" resultid="7428" />
                    <RANKING order="4" place="4" resultid="8679" />
                    <RANKING order="5" place="5" resultid="9465" />
                    <RANKING order="6" place="-1" resultid="9466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1671" agemax="239" agemin="200" name="Kat D 200-239">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9644" />
                    <RANKING order="2" place="2" resultid="7426" />
                    <RANKING order="3" place="3" resultid="6515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1672" agemax="279" agemin="240" name="Kat E 240-279">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8994" />
                    <RANKING order="2" place="2" resultid="8805" />
                    <RANKING order="3" place="3" resultid="6704" />
                    <RANKING order="4" place="4" resultid="7424" />
                    <RANKING order="5" place="5" resultid="3318" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1673" agemax="-1" agemin="280" name="Kat F 280 +">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8804" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10927" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10928" daytime="10:53" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10929" daytime="10:57" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1674" daytime="11:00" gender="F" number="39" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2795" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2796" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3228" />
                    <RANKING order="2" place="2" resultid="3515" />
                    <RANKING order="3" place="-1" resultid="3637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2797" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8379" />
                    <RANKING order="2" place="2" resultid="9864" />
                    <RANKING order="3" place="3" resultid="8551" />
                    <RANKING order="4" place="4" resultid="8486" />
                    <RANKING order="5" place="5" resultid="8586" />
                    <RANKING order="6" place="6" resultid="6446" />
                    <RANKING order="7" place="-1" resultid="7373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2798" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6341" />
                    <RANKING order="2" place="2" resultid="8643" />
                    <RANKING order="3" place="3" resultid="6501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2799" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8831" />
                    <RANKING order="2" place="2" resultid="7906" />
                    <RANKING order="3" place="3" resultid="8496" />
                    <RANKING order="4" place="4" resultid="9364" />
                    <RANKING order="5" place="5" resultid="3289" />
                    <RANKING order="6" place="6" resultid="6768" />
                    <RANKING order="7" place="-1" resultid="8309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2800" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7360" />
                    <RANKING order="2" place="2" resultid="9373" />
                    <RANKING order="3" place="3" resultid="7572" />
                    <RANKING order="4" place="-1" resultid="3240" />
                    <RANKING order="5" place="-1" resultid="8793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2801" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9124" />
                    <RANKING order="2" place="2" resultid="6415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2802" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7353" />
                    <RANKING order="2" place="2" resultid="8092" />
                    <RANKING order="3" place="3" resultid="8935" />
                    <RANKING order="4" place="4" resultid="6453" />
                    <RANKING order="5" place="-1" resultid="6669" />
                    <RANKING order="6" place="-1" resultid="8944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2803" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7346" />
                    <RANKING order="2" place="2" resultid="6688" />
                    <RANKING order="3" place="3" resultid="3208" />
                    <RANKING order="4" place="4" resultid="9609" />
                    <RANKING order="5" place="5" resultid="6460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2804" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4583" />
                    <RANKING order="2" place="2" resultid="8572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2805" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8770" />
                    <RANKING order="2" place="2" resultid="7984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2806" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2807" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2808" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2809" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2810" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10930" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10931" daytime="11:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10932" daytime="11:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10933" daytime="11:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10934" daytime="11:38" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1623" daytime="10:21" gender="F" number="36" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2763" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9388" />
                    <RANKING order="2" place="2" resultid="10130" />
                    <RANKING order="3" place="3" resultid="9492" />
                    <RANKING order="4" place="4" resultid="3312" />
                    <RANKING order="5" place="5" resultid="3199" />
                    <RANKING order="6" place="6" resultid="7091" />
                    <RANKING order="7" place="7" resultid="9440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2764" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2765" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6787" />
                    <RANKING order="2" place="2" resultid="7938" />
                    <RANKING order="3" place="3" resultid="9847" />
                    <RANKING order="4" place="4" resultid="10296" />
                    <RANKING order="5" place="5" resultid="8378" />
                    <RANKING order="6" place="6" resultid="8613" />
                    <RANKING order="7" place="7" resultid="8917" />
                    <RANKING order="8" place="8" resultid="8847" />
                    <RANKING order="9" place="9" resultid="9873" />
                    <RANKING order="10" place="10" resultid="8664" />
                    <RANKING order="11" place="11" resultid="3848" />
                    <RANKING order="12" place="12" resultid="9855" />
                    <RANKING order="13" place="-1" resultid="6594" />
                    <RANKING order="14" place="-1" resultid="8485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2766" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7968" />
                    <RANKING order="2" place="2" resultid="6327" />
                    <RANKING order="3" place="3" resultid="8271" />
                    <RANKING order="4" place="4" resultid="7368" />
                    <RANKING order="5" place="5" resultid="8028" />
                    <RANKING order="6" place="6" resultid="8855" />
                    <RANKING order="7" place="7" resultid="6500" />
                    <RANKING order="8" place="-1" resultid="9393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2767" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6319" />
                    <RANKING order="2" place="2" resultid="9489" />
                    <RANKING order="3" place="3" resultid="9535" />
                    <RANKING order="4" place="4" resultid="9414" />
                    <RANKING order="5" place="5" resultid="6585" />
                    <RANKING order="6" place="6" resultid="7835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2768" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3649" />
                    <RANKING order="2" place="2" resultid="8792" />
                    <RANKING order="3" place="3" resultid="8627" />
                    <RANKING order="4" place="4" resultid="10108" />
                    <RANKING order="5" place="5" resultid="3269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2769" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6609" />
                    <RANKING order="2" place="2" resultid="8075" />
                    <RANKING order="3" place="3" resultid="6414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2770" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8943" />
                    <RANKING order="2" place="2" resultid="9356" />
                    <RANKING order="3" place="3" resultid="6488" />
                    <RANKING order="4" place="4" resultid="6495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2771" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9581" />
                    <RANKING order="2" place="2" resultid="7338" />
                    <RANKING order="3" place="3" resultid="10096" />
                    <RANKING order="4" place="4" resultid="8313" />
                    <RANKING order="5" place="5" resultid="7349" />
                    <RANKING order="6" place="6" resultid="10609" />
                    <RANKING order="7" place="-1" resultid="7564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2772" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4582" />
                    <RANKING order="2" place="2" resultid="7482" />
                    <RANKING order="3" place="3" resultid="9071" />
                    <RANKING order="4" place="-1" resultid="7327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2773" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8764" />
                    <RANKING order="2" place="2" resultid="6629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2774" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2775" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2776" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2777" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2778" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10905" daytime="10:21" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10906" daytime="10:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10907" daytime="10:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10908" daytime="10:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10909" daytime="10:27" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10910" daytime="10:28" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10911" daytime="10:29" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1578" daytime="09:09" gender="M" number="33" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2715" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10316" />
                    <RANKING order="2" place="2" resultid="7087" />
                    <RANKING order="3" place="3" resultid="8420" />
                    <RANKING order="4" place="4" resultid="7600" />
                    <RANKING order="5" place="-1" resultid="7149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2716" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7594" />
                    <RANKING order="2" place="2" resultid="8472" />
                    <RANKING order="3" place="3" resultid="7066" />
                    <RANKING order="4" place="4" resultid="7135" />
                    <RANKING order="5" place="-1" resultid="6853" />
                    <RANKING order="6" place="-1" resultid="7743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2717" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6561" />
                    <RANKING order="2" place="2" resultid="8838" />
                    <RANKING order="3" place="3" resultid="3881" />
                    <RANKING order="4" place="4" resultid="9801" />
                    <RANKING order="5" place="5" resultid="6885" />
                    <RANKING order="6" place="6" resultid="7631" />
                    <RANKING order="7" place="-1" resultid="6804" />
                    <RANKING order="8" place="-1" resultid="6962" />
                    <RANKING order="9" place="-1" resultid="8971" />
                    <RANKING order="10" place="-1" resultid="9900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2718" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9886" />
                    <RANKING order="2" place="2" resultid="9589" />
                    <RANKING order="3" place="3" resultid="6399" />
                    <RANKING order="4" place="4" resultid="8910" />
                    <RANKING order="5" place="5" resultid="6872" />
                    <RANKING order="6" place="6" resultid="8844" />
                    <RANKING order="7" place="7" resultid="8529" />
                    <RANKING order="8" place="8" resultid="3254" />
                    <RANKING order="9" place="-1" resultid="8366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2719" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6780" />
                    <RANKING order="2" place="2" resultid="8081" />
                    <RANKING order="3" place="3" resultid="8025" />
                    <RANKING order="4" place="4" resultid="10276" />
                    <RANKING order="5" place="5" resultid="10258" />
                    <RANKING order="6" place="-1" resultid="7648" />
                    <RANKING order="7" place="-1" resultid="8262" />
                    <RANKING order="8" place="-1" resultid="8453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2720" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8204" />
                    <RANKING order="2" place="2" resultid="7785" />
                    <RANKING order="3" place="3" resultid="6986" />
                    <RANKING order="4" place="4" resultid="10170" />
                    <RANKING order="5" place="5" resultid="8236" />
                    <RANKING order="6" place="6" resultid="8208" />
                    <RANKING order="7" place="-1" resultid="6975" />
                    <RANKING order="8" place="-1" resultid="8301" />
                    <RANKING order="9" place="-1" resultid="8429" />
                    <RANKING order="10" place="-1" resultid="8650" />
                    <RANKING order="11" place="-1" resultid="9785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2721" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6432" />
                    <RANKING order="2" place="2" resultid="3659" />
                    <RANKING order="3" place="3" resultid="6440" />
                    <RANKING order="4" place="4" resultid="10581" />
                    <RANKING order="5" place="5" resultid="7588" />
                    <RANKING order="6" place="6" resultid="9453" />
                    <RANKING order="7" place="7" resultid="8501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2722" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7620" />
                    <RANKING order="2" place="2" resultid="6694" />
                    <RANKING order="3" place="3" resultid="8516" />
                    <RANKING order="4" place="4" resultid="6352" />
                    <RANKING order="5" place="-1" resultid="8049" />
                    <RANKING order="6" place="-1" resultid="9110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2723" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8987" />
                    <RANKING order="2" place="2" resultid="7927" />
                    <RANKING order="3" place="3" resultid="6774" />
                    <RANKING order="4" place="4" resultid="6310" />
                    <RANKING order="5" place="5" resultid="6755" />
                    <RANKING order="6" place="6" resultid="8901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2724" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8336" />
                    <RANKING order="2" place="2" resultid="9841" />
                    <RANKING order="3" place="3" resultid="8359" />
                    <RANKING order="4" place="-1" resultid="6532" />
                    <RANKING order="5" place="-1" resultid="7558" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2725" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8927" />
                    <RANKING order="2" place="2" resultid="7778" />
                    <RANKING order="3" place="3" resultid="6620" />
                    <RANKING order="4" place="-1" resultid="7991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2726" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6375" />
                    <RANKING order="2" place="2" resultid="7977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2727" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2728" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2729" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2730" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10885" daytime="09:09" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10886" daytime="09:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10887" daytime="09:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10888" daytime="09:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10889" daytime="09:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10890" daytime="09:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10891" daytime="09:21" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10892" daytime="09:23" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1593" daytime="09:25" gender="F" number="34" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2731" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9640" />
                    <RANKING order="2" place="2" resultid="9637" />
                    <RANKING order="3" place="3" resultid="10557" />
                    <RANKING order="4" place="4" resultid="10129" />
                    <RANKING order="5" place="5" resultid="3198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2732" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7762" />
                    <RANKING order="2" place="2" resultid="3210" />
                    <RANKING order="3" place="3" resultid="3514" />
                    <RANKING order="4" place="-1" resultid="3636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2733" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9863" />
                    <RANKING order="2" place="2" resultid="9854" />
                    <RANKING order="3" place="3" resultid="8585" />
                    <RANKING order="4" place="-1" resultid="9349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2734" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3870" />
                    <RANKING order="2" place="2" resultid="7662" />
                    <RANKING order="3" place="3" resultid="8854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2735" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8957" />
                    <RANKING order="2" place="2" resultid="8830" />
                    <RANKING order="3" place="3" resultid="7160" />
                    <RANKING order="4" place="4" resultid="6589" />
                    <RANKING order="5" place="5" resultid="7658" />
                    <RANKING order="6" place="6" resultid="8308" />
                    <RANKING order="7" place="7" resultid="9363" />
                    <RANKING order="8" place="8" resultid="9655" />
                    <RANKING order="9" place="-1" resultid="3262" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2736" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7359" />
                    <RANKING order="2" place="2" resultid="6679" />
                    <RANKING order="3" place="3" resultid="3268" />
                    <RANKING order="4" place="4" resultid="7571" />
                    <RANKING order="5" place="-1" resultid="6751" />
                    <RANKING order="6" place="-1" resultid="8965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2737" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9123" />
                    <RANKING order="2" place="2" resultid="6361" />
                    <RANKING order="3" place="3" resultid="6293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2738" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8091" />
                    <RANKING order="2" place="2" resultid="9114" />
                    <RANKING order="3" place="3" resultid="6487" />
                    <RANKING order="4" place="4" resultid="9600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2739" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7345" />
                    <RANKING order="2" place="2" resultid="3219" />
                    <RANKING order="3" place="3" resultid="6459" />
                    <RANKING order="4" place="4" resultid="9608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2740" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2741" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2742" agemax="79" agemin="75" name="Kat K 75-79" />
                <AGEGROUP agegroupid="2743" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2744" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2745" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2746" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10893" daytime="09:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10894" daytime="09:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10895" daytime="09:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10896" daytime="09:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10897" daytime="09:45" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1695" daytime="11:45" gender="M" number="40" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2811" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9522" />
                    <RANKING order="2" place="2" resultid="10651" />
                    <RANKING order="3" place="3" resultid="7088" />
                    <RANKING order="4" place="4" resultid="6479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2812" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3644" />
                    <RANKING order="2" place="2" resultid="7067" />
                    <RANKING order="3" place="3" resultid="7595" />
                    <RANKING order="4" place="4" resultid="7744" />
                    <RANKING order="5" place="5" resultid="3843" />
                    <RANKING order="6" place="-1" resultid="6864" />
                    <RANKING order="7" place="-1" resultid="7075" />
                    <RANKING order="8" place="-1" resultid="7769" />
                    <RANKING order="9" place="-1" resultid="8224" />
                    <RANKING order="10" place="-1" resultid="9915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2813" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7155" />
                    <RANKING order="2" place="2" resultid="9105" />
                    <RANKING order="3" place="3" resultid="8555" />
                    <RANKING order="4" place="4" resultid="8372" />
                    <RANKING order="5" place="5" resultid="6805" />
                    <RANKING order="6" place="6" resultid="8592" />
                    <RANKING order="7" place="7" resultid="3882" />
                    <RANKING order="8" place="8" resultid="9530" />
                    <RANKING order="9" place="9" resultid="3893" />
                    <RANKING order="10" place="10" resultid="6060" />
                    <RANKING order="11" place="-1" resultid="6562" />
                    <RANKING order="12" place="-1" resultid="8839" />
                    <RANKING order="13" place="-1" resultid="10261" />
                    <RANKING order="14" place="-1" resultid="10953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2814" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9590" />
                    <RANKING order="2" place="2" resultid="8447" />
                    <RANKING order="3" place="3" resultid="8576" />
                    <RANKING order="4" place="4" resultid="6891" />
                    <RANKING order="5" place="5" resultid="7641" />
                    <RANKING order="6" place="6" resultid="8530" />
                    <RANKING order="7" place="7" resultid="6513" />
                    <RANKING order="8" place="8" resultid="8609" />
                    <RANKING order="9" place="9" resultid="10041" />
                    <RANKING order="10" place="10" resultid="10664" />
                    <RANKING order="11" place="-1" resultid="8344" />
                    <RANKING order="12" place="-1" resultid="8367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2815" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8082" />
                    <RANKING order="2" place="2" resultid="7649" />
                    <RANKING order="3" place="3" resultid="6812" />
                    <RANKING order="4" place="4" resultid="9101" />
                    <RANKING order="5" place="5" resultid="6575" />
                    <RANKING order="6" place="6" resultid="8245" />
                    <RANKING order="7" place="7" resultid="7158" />
                    <RANKING order="8" place="8" resultid="7829" />
                    <RANKING order="9" place="9" resultid="8494" />
                    <RANKING order="10" place="10" resultid="3860" />
                    <RANKING order="11" place="11" resultid="7675" />
                    <RANKING order="12" place="12" resultid="7003" />
                    <RANKING order="13" place="13" resultid="3185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2816" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7413" />
                    <RANKING order="2" place="2" resultid="3299" />
                    <RANKING order="3" place="3" resultid="8430" />
                    <RANKING order="4" place="4" resultid="4574" />
                    <RANKING order="5" place="5" resultid="9786" />
                    <RANKING order="6" place="6" resultid="7625" />
                    <RANKING order="7" place="7" resultid="8481" />
                    <RANKING order="8" place="-1" resultid="6425" />
                    <RANKING order="9" place="-1" resultid="8205" />
                    <RANKING order="10" place="-1" resultid="8302" />
                    <RANKING order="11" place="-1" resultid="9817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2817" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6433" />
                    <RANKING order="2" place="2" resultid="7589" />
                    <RANKING order="3" place="3" resultid="7408" />
                    <RANKING order="4" place="4" resultid="8538" />
                    <RANKING order="5" place="5" resultid="7609" />
                    <RANKING order="6" place="6" resultid="7401" />
                    <RANKING order="7" place="7" resultid="9812" />
                    <RANKING order="8" place="-1" resultid="6347" />
                    <RANKING order="9" place="-1" resultid="8322" />
                    <RANKING order="10" place="-1" resultid="9454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2818" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8509" />
                    <RANKING order="2" place="2" resultid="9622" />
                    <RANKING order="3" place="3" resultid="7621" />
                    <RANKING order="4" place="4" resultid="6408" />
                    <RANKING order="5" place="5" resultid="8517" />
                    <RANKING order="6" place="6" resultid="7943" />
                    <RANKING order="7" place="-1" resultid="7580" />
                    <RANKING order="8" place="-1" resultid="8050" />
                    <RANKING order="9" place="-1" resultid="9119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2819" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8988" />
                    <RANKING order="2" place="2" resultid="7389" />
                    <RANKING order="3" place="3" resultid="10271" />
                    <RANKING order="4" place="4" resultid="6795" />
                    <RANKING order="5" place="5" resultid="4565" />
                    <RANKING order="6" place="6" resultid="8097" />
                    <RANKING order="7" place="7" resultid="8630" />
                    <RANKING order="8" place="8" resultid="8902" />
                    <RANKING order="9" place="9" resultid="8889" />
                    <RANKING order="10" place="-1" resultid="6385" />
                    <RANKING order="11" place="-1" resultid="7531" />
                    <RANKING order="12" place="-1" resultid="8000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2820" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8068" />
                    <RANKING order="2" place="2" resultid="8949" />
                    <RANKING order="3" place="3" resultid="7554" />
                    <RANKING order="4" place="4" resultid="9037" />
                    <RANKING order="5" place="5" resultid="9842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2821" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6621" />
                    <RANKING order="2" place="2" resultid="8584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2822" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8767" />
                    <RANKING order="2" place="2" resultid="6647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2823" agemax="84" agemin="80" name="Kat L 80-84" />
                <AGEGROUP agegroupid="2824" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2825" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2826" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10935" daytime="11:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10936" daytime="11:57" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10937" daytime="12:09" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10938" daytime="12:17" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10939" daytime="12:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10940" daytime="12:31" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10941" daytime="12:37" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10942" daytime="12:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10943" daytime="12:49" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10944" daytime="12:55" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10945" daytime="13:01" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1638" daytime="10:31" gender="M" number="37" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2779" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6847" />
                    <RANKING order="2" place="2" resultid="9523" />
                    <RANKING order="3" place="3" resultid="6478" />
                    <RANKING order="4" place="4" resultid="10317" />
                    <RANKING order="5" place="5" resultid="10120" />
                    <RANKING order="6" place="6" resultid="8421" />
                    <RANKING order="7" place="7" resultid="9834" />
                    <RANKING order="8" place="8" resultid="10234" />
                    <RANKING order="9" place="-1" resultid="7150" />
                    <RANKING order="10" place="-1" resultid="10310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2780" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6817" />
                    <RANKING order="2" place="2" resultid="7009" />
                    <RANKING order="3" place="3" resultid="7074" />
                    <RANKING order="4" place="4" resultid="6301" />
                    <RANKING order="5" place="5" resultid="3525" />
                    <RANKING order="6" place="6" resultid="7140" />
                    <RANKING order="7" place="7" resultid="3842" />
                    <RANKING order="8" place="8" resultid="9402" />
                    <RANKING order="9" place="9" resultid="9418" />
                    <RANKING order="10" place="-1" resultid="8473" />
                    <RANKING order="11" place="-1" resultid="6858" />
                    <RANKING order="12" place="-1" resultid="8223" />
                    <RANKING order="13" place="-1" resultid="10567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2781" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8605" />
                    <RANKING order="2" place="2" resultid="9878" />
                    <RANKING order="3" place="3" resultid="7095" />
                    <RANKING order="4" place="4" resultid="7793" />
                    <RANKING order="5" place="5" resultid="6907" />
                    <RANKING order="6" place="6" resultid="6304" />
                    <RANKING order="7" place="7" resultid="3829" />
                    <RANKING order="8" place="8" resultid="7632" />
                    <RANKING order="9" place="9" resultid="8863" />
                    <RANKING order="10" place="10" resultid="9802" />
                    <RANKING order="11" place="11" resultid="9822" />
                    <RANKING order="12" place="-1" resultid="6963" />
                    <RANKING order="13" place="-1" resultid="8972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2782" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8911" />
                    <RANKING order="2" place="2" resultid="8562" />
                    <RANKING order="3" place="3" resultid="9617" />
                    <RANKING order="4" place="4" resultid="6877" />
                    <RANKING order="5" place="5" resultid="10563" />
                    <RANKING order="6" place="6" resultid="6901" />
                    <RANKING order="7" place="7" resultid="6918" />
                    <RANKING order="8" place="8" resultid="7002" />
                    <RANKING order="9" place="9" resultid="7651" />
                    <RANKING order="10" place="10" resultid="10040" />
                    <RANKING order="11" place="11" resultid="6999" />
                    <RANKING order="12" place="12" resultid="10663" />
                    <RANKING order="13" place="13" resultid="3255" />
                    <RANKING order="14" place="-1" resultid="10291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2783" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8263" />
                    <RANKING order="2" place="2" resultid="8568" />
                    <RANKING order="3" place="3" resultid="8250" />
                    <RANKING order="4" place="4" resultid="8596" />
                    <RANKING order="5" place="5" resultid="8059" />
                    <RANKING order="6" place="6" resultid="6612" />
                    <RANKING order="7" place="7" resultid="6580" />
                    <RANKING order="8" place="8" resultid="3184" />
                    <RANKING order="9" place="9" resultid="10259" />
                    <RANKING order="10" place="10" resultid="3859" />
                    <RANKING order="11" place="11" resultid="8493" />
                    <RANKING order="12" place="12" resultid="8020" />
                    <RANKING order="13" place="13" resultid="8015" />
                    <RANKING order="14" place="14" resultid="9793" />
                    <RANKING order="15" place="-1" resultid="6971" />
                    <RANKING order="16" place="-1" resultid="7798" />
                    <RANKING order="17" place="-1" resultid="8010" />
                    <RANKING order="18" place="-1" resultid="8454" />
                    <RANKING order="19" place="-1" resultid="10161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2784" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7786" />
                    <RANKING order="2" place="2" resultid="6981" />
                    <RANKING order="3" place="3" resultid="8231" />
                    <RANKING order="4" place="4" resultid="3298" />
                    <RANKING order="5" place="5" resultid="8237" />
                    <RANKING order="6" place="6" resultid="8256" />
                    <RANKING order="7" place="7" resultid="7789" />
                    <RANKING order="8" place="8" resultid="6745" />
                    <RANKING order="9" place="9" resultid="8480" />
                    <RANKING order="10" place="10" resultid="9409" />
                    <RANKING order="11" place="-1" resultid="7025" />
                    <RANKING order="12" place="-1" resultid="3888" />
                    <RANKING order="13" place="-1" resultid="6424" />
                    <RANKING order="14" place="-1" resultid="6976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2785" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6287" />
                    <RANKING order="2" place="2" resultid="7407" />
                    <RANKING order="3" place="3" resultid="6535" />
                    <RANKING order="4" place="4" resultid="6808" />
                    <RANKING order="5" place="5" resultid="10582" />
                    <RANKING order="6" place="6" resultid="7400" />
                    <RANKING order="7" place="7" resultid="6634" />
                    <RANKING order="8" place="8" resultid="8502" />
                    <RANKING order="9" place="9" resultid="9789" />
                    <RANKING order="10" place="10" resultid="9811" />
                    <RANKING order="11" place="-1" resultid="6441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2786" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6538" />
                    <RANKING order="2" place="2" resultid="9921" />
                    <RANKING order="3" place="3" resultid="6695" />
                    <RANKING order="4" place="4" resultid="9627" />
                    <RANKING order="5" place="5" resultid="9111" />
                    <RANKING order="6" place="6" resultid="8921" />
                    <RANKING order="7" place="7" resultid="7393" />
                    <RANKING order="8" place="8" resultid="8953" />
                    <RANKING order="9" place="9" resultid="6353" />
                    <RANKING order="10" place="-1" resultid="7548" />
                    <RANKING order="11" place="-1" resultid="8508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2787" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10575" />
                    <RANKING order="2" place="2" resultid="10332" />
                    <RANKING order="3" place="3" resultid="7928" />
                    <RANKING order="4" place="4" resultid="9075" />
                    <RANKING order="5" place="5" resultid="6311" />
                    <RANKING order="6" place="6" resultid="9127" />
                    <RANKING order="7" place="7" resultid="7388" />
                    <RANKING order="8" place="8" resultid="6555" />
                    <RANKING order="9" place="-1" resultid="6384" />
                    <RANKING order="10" place="-1" resultid="8096" />
                    <RANKING order="11" place="-1" resultid="10270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2788" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8635" />
                    <RANKING order="2" place="2" resultid="8893" />
                    <RANKING order="3" place="3" resultid="8948" />
                    <RANKING order="4" place="4" resultid="7381" />
                    <RANKING order="5" place="5" resultid="8993" />
                    <RANKING order="6" place="6" resultid="8384" />
                    <RANKING order="7" place="7" resultid="3233" />
                    <RANKING order="8" place="-1" resultid="7559" />
                    <RANKING order="9" place="-1" resultid="7915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2789" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7480" />
                    <RANKING order="2" place="2" resultid="7779" />
                    <RANKING order="3" place="3" resultid="7377" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2790" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6376" />
                    <RANKING order="2" place="2" resultid="8759" />
                    <RANKING order="3" place="3" resultid="9066" />
                    <RANKING order="4" place="4" resultid="8435" />
                    <RANKING order="5" place="5" resultid="8211" />
                    <RANKING order="6" place="6" resultid="8319" />
                    <RANKING order="7" place="7" resultid="6646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2791" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9080" />
                    <RANKING order="2" place="2" resultid="8353" />
                    <RANKING order="3" place="-1" resultid="7755" />
                    <RANKING order="4" place="-1" resultid="8546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2792" agemax="89" agemin="85" name="Kat M  85-89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3248" />
                    <RANKING order="2" place="2" resultid="3164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2793" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2794" agemax="99" agemin="95" name="Kat O 95-99">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8884" />
                    <RANKING order="2" place="-1" resultid="7325" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10912" daytime="10:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10913" daytime="10:33" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10914" daytime="10:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10915" daytime="10:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10916" daytime="10:37" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10917" daytime="10:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10918" daytime="10:39" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10919" daytime="10:41" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10920" daytime="10:42" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10921" daytime="10:43" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10922" daytime="10:44" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10923" daytime="10:45" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="10924" daytime="10:46" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="10925" daytime="10:47" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="10926" daytime="10:48" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1608" daytime="09:49" gender="M" number="35" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2747" agemax="24" agemin="20" name="Kat 0 - 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10650" />
                    <RANKING order="2" place="2" resultid="9833" />
                    <RANKING order="3" place="3" resultid="10119" />
                    <RANKING order="4" place="-1" resultid="10309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2748" agemax="29" agemin="25" name="Kat A - 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7073" />
                    <RANKING order="2" place="2" resultid="3524" />
                    <RANKING order="3" place="-1" resultid="9914" />
                    <RANKING order="4" place="-1" resultid="10091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2749" agemax="34" agemin="30" name="Kat B - 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6603" />
                    <RANKING order="2" place="2" resultid="6897" />
                    <RANKING order="3" place="3" resultid="9895" />
                    <RANKING order="4" place="4" resultid="10952" />
                    <RANKING order="5" place="5" resultid="8862" />
                    <RANKING order="6" place="6" resultid="6059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2750" agemax="39" agemin="35" name="Kat C 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9887" />
                    <RANKING order="2" place="2" resultid="8655" />
                    <RANKING order="3" place="3" resultid="9632" />
                    <RANKING order="4" place="4" resultid="8978" />
                    <RANKING order="5" place="5" resultid="8446" />
                    <RANKING order="6" place="6" resultid="9431" />
                    <RANKING order="7" place="7" resultid="8343" />
                    <RANKING order="8" place="8" resultid="6917" />
                    <RANKING order="9" place="-1" resultid="8330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2751" agemax="44" agemin="40" name="Kat D 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10241" />
                    <RANKING order="2" place="2" resultid="9514" />
                    <RANKING order="3" place="3" resultid="9100" />
                    <RANKING order="4" place="4" resultid="8058" />
                    <RANKING order="5" place="5" resultid="6574" />
                    <RANKING order="6" place="6" resultid="8244" />
                    <RANKING order="7" place="-1" resultid="7674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2752" agemax="49" agemin="45" name="Kat E 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8201" />
                    <RANKING order="2" place="2" resultid="3790" />
                    <RANKING order="3" place="3" resultid="7417" />
                    <RANKING order="4" place="4" resultid="6744" />
                    <RANKING order="5" place="5" resultid="4573" />
                    <RANKING order="6" place="-1" resultid="6994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2753" agemax="54" agemin="50" name="Kat F 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10166" />
                    <RANKING order="2" place="2" resultid="8524" />
                    <RANKING order="3" place="3" resultid="6346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2754" agemax="59" agemin="55" name="Kat G 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7748" />
                    <RANKING order="2" place="2" resultid="9920" />
                    <RANKING order="3" place="3" resultid="6764" />
                    <RANKING order="4" place="4" resultid="8778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2755" agemax="64" agemin="60" name="Kat H 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8535" />
                    <RANKING order="2" place="2" resultid="4564" />
                    <RANKING order="3" place="3" resultid="7999" />
                    <RANKING order="4" place="4" resultid="6794" />
                    <RANKING order="5" place="5" resultid="7530" />
                    <RANKING order="6" place="6" resultid="6507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2756" agemax="69" agemin="65" name="Kat I 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8461" />
                    <RANKING order="2" place="2" resultid="8067" />
                    <RANKING order="3" place="3" resultid="9036" />
                    <RANKING order="4" place="4" resultid="3282" />
                    <RANKING order="5" place="5" resultid="8360" />
                    <RANKING order="6" place="-1" resultid="6533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2757" agemax="74" agemin="70" name="Kat J 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7832" />
                    <RANKING order="2" place="2" resultid="8797" />
                    <RANKING order="3" place="-1" resultid="7992" />
                    <RANKING order="4" place="-1" resultid="8583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2758" agemax="79" agemin="75" name="Kat K 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7978" />
                    <RANKING order="2" place="2" resultid="8318" />
                    <RANKING order="3" place="3" resultid="8349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2759" agemax="84" agemin="80" name="Kat L 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7754" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2760" agemax="89" agemin="85" name="Kat M  85-89" />
                <AGEGROUP agegroupid="2761" agemax="94" agemin="90" name="Kat N  90-94" />
                <AGEGROUP agegroupid="2762" agemax="99" agemin="95" name="Kat O 95-99" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10898" daytime="09:49" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10899" daytime="09:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10900" daytime="10:01" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10901" daytime="10:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10902" daytime="10:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10903" daytime="10:14" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10904" daytime="10:17" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="ALTEM" nation="RUS" clubid="11097" name="Alex Fitness ">
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Timur" gender="M" lastname="Podmarev" nation="POL" athleteid="6225">
              <RESULTS>
                <RESULT eventid="1190" points="386" swimtime="00:02:36.57" resultid="10571" heatid="10727" lane="4" entrytime="00:02:37.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:15.44" />
                    <SPLIT distance="150" swimtime="00:01:57.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="442" swimtime="00:02:46.71" resultid="10572" heatid="10763" lane="3" entrytime="00:02:45.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="100" swimtime="00:01:20.14" />
                    <SPLIT distance="150" swimtime="00:02:03.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="326" swimtime="00:02:41.88" resultid="10573" heatid="10795" lane="5" entrytime="00:02:40.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:16.34" />
                    <SPLIT distance="150" swimtime="00:01:59.95" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Europy Masters  Mężczyzn w  kat H 60-64  lata" eventid="1392" points="424" swimtime="00:01:15.99" resultid="10574" heatid="10818" lane="2" entrytime="00:01:14.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="469" swimtime="00:00:34.00" resultid="10575" heatid="10924" lane="6" entrytime="00:00:33.87" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AQKYI" nation="UKR" clubid="4945" name="Aqua Masters Kyiv">
          <CONTACT city="Kyiv" email="romaniokiev@gmail.com" name="Rallo Oleksandr" phone="+38 050 3535704" zip="03000" />
          <ATHLETES>
            <ATHLETE birthdate="1957-10-08" firstname="Volodymyr" gender="M" lastname="Turchyn" nation="UKR" athleteid="4946">
              <RESULTS>
                <RESULT eventid="1160" points="274" swimtime="00:00:32.16" resultid="6771" heatid="10699" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="6772" heatid="10778" lane="9" entrytime="00:01:12.00" />
                <RESULT eventid="1422" points="304" swimtime="00:00:33.33" resultid="6773" heatid="10831" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1578" points="151" swimtime="00:01:33.36" resultid="6774" heatid="10887" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AQOLS" nation="POL" region="WAR" clubid="5020" name="Aquasfera Masters Olsztyn">
          <CONTACT email="annamariaaneczka@gmail.com" name="Goździejewska Anna" />
          <ATHLETES>
            <ATHLETE birthdate="1992-02-28" firstname="Maciej" gender="M" lastname="Zembrzuski" nation="POL" athleteid="5055">
              <RESULTS>
                <RESULT eventid="1160" points="627" swimtime="00:00:24.42" resultid="7590" heatid="10710" lane="8" entrytime="00:00:25.49" />
                <RESULT eventid="1302" points="651" swimtime="00:00:54.11" resultid="7591" heatid="10788" lane="3" entrytime="00:00:54.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="632" swimtime="00:00:26.13" resultid="7592" heatid="10838" lane="0" entrytime="00:00:26.30" />
                <RESULT eventid="1482" points="559" swimtime="00:02:03.82" resultid="7593" heatid="10866" lane="5" entrytime="00:01:59.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                    <SPLIT distance="100" swimtime="00:00:59.90" />
                    <SPLIT distance="150" swimtime="00:01:32.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="595" swimtime="00:00:59.21" resultid="7594" heatid="10892" lane="5" entrytime="00:00:58.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="449" swimtime="00:04:47.23" resultid="7595" heatid="10945" lane="6" entrytime="00:04:32.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:01:05.04" />
                    <SPLIT distance="150" swimtime="00:01:40.13" />
                    <SPLIT distance="200" swimtime="00:02:15.70" />
                    <SPLIT distance="250" swimtime="00:02:51.97" />
                    <SPLIT distance="300" swimtime="00:03:29.89" />
                    <SPLIT distance="350" swimtime="00:04:09.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-26" firstname="Grzegorz" gender="M" lastname="Kalinowski" nation="POL" athleteid="5106">
              <RESULTS>
                <RESULT eventid="1160" points="311" swimtime="00:00:30.85" resultid="7633" heatid="10699" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1242" points="238" swimtime="00:00:38.75" resultid="7634" heatid="10747" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1302" points="308" swimtime="00:01:09.46" resultid="7635" heatid="10779" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="220" swimtime="00:01:25.78" resultid="7636" heatid="10846" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-10-01" firstname="Katarzyna" gender="F" lastname="Klajbor" nation="POL" athleteid="5035">
              <RESULTS>
                <RESULT eventid="1059" points="293" swimtime="00:12:09.44" resultid="7573" heatid="10667" lane="0" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                    <SPLIT distance="100" swimtime="00:01:25.35" />
                    <SPLIT distance="150" swimtime="00:02:11.12" />
                    <SPLIT distance="200" swimtime="00:02:56.56" />
                    <SPLIT distance="250" swimtime="00:03:42.93" />
                    <SPLIT distance="300" swimtime="00:04:28.75" />
                    <SPLIT distance="350" swimtime="00:05:14.49" />
                    <SPLIT distance="400" swimtime="00:06:00.62" />
                    <SPLIT distance="450" swimtime="00:06:47.38" />
                    <SPLIT distance="500" swimtime="00:07:33.81" />
                    <SPLIT distance="550" swimtime="00:08:20.39" />
                    <SPLIT distance="600" swimtime="00:09:07.06" />
                    <SPLIT distance="650" swimtime="00:09:53.35" />
                    <SPLIT distance="700" swimtime="00:10:39.76" />
                    <SPLIT distance="750" swimtime="00:11:25.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="287" swimtime="00:01:18.88" resultid="7574" heatid="10766" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-08-31" firstname="Iwona" gender="F" lastname="Bardzicka" nation="POL" athleteid="5021">
              <RESULTS>
                <RESULT eventid="1059" points="56" swimtime="00:21:01.14" resultid="7561" heatid="10666" lane="9" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.35" />
                    <SPLIT distance="100" swimtime="00:02:25.42" />
                    <SPLIT distance="150" swimtime="00:03:40.90" />
                    <SPLIT distance="200" swimtime="00:04:57.87" />
                    <SPLIT distance="250" swimtime="00:06:16.00" />
                    <SPLIT distance="300" swimtime="00:07:35.06" />
                    <SPLIT distance="350" swimtime="00:08:53.91" />
                    <SPLIT distance="400" swimtime="00:10:14.04" />
                    <SPLIT distance="450" swimtime="00:11:35.10" />
                    <SPLIT distance="500" swimtime="00:12:56.07" />
                    <SPLIT distance="550" swimtime="00:14:17.75" />
                    <SPLIT distance="600" swimtime="00:15:39.35" />
                    <SPLIT distance="650" swimtime="00:17:01.41" />
                    <SPLIT distance="700" swimtime="00:18:23.36" />
                    <SPLIT distance="750" swimtime="00:19:43.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="108" swimtime="00:04:51.96" resultid="7562" heatid="10753" lane="1" entrytime="00:04:42.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.80" />
                    <SPLIT distance="100" swimtime="00:02:18.07" />
                    <SPLIT distance="150" swimtime="00:03:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="111" swimtime="00:02:13.59" resultid="7563" heatid="10804" lane="9" entrytime="00:02:09.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="7564" heatid="10906" lane="6" entrytime="00:00:58.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-03-18" firstname="Danuta" gender="F" lastname="Wegen" nation="POL" athleteid="5026">
              <RESULTS>
                <RESULT eventid="1059" points="90" swimtime="00:17:58.30" resultid="7565" heatid="10666" lane="5" entrytime="00:15:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.94" />
                    <SPLIT distance="100" swimtime="00:01:58.64" />
                    <SPLIT distance="150" swimtime="00:03:07.33" />
                    <SPLIT distance="200" swimtime="00:04:16.61" />
                    <SPLIT distance="250" swimtime="00:05:25.95" />
                    <SPLIT distance="300" swimtime="00:06:34.70" />
                    <SPLIT distance="350" swimtime="00:07:43.35" />
                    <SPLIT distance="400" swimtime="00:08:51.85" />
                    <SPLIT distance="450" swimtime="00:10:02.21" />
                    <SPLIT distance="500" swimtime="00:11:10.61" />
                    <SPLIT distance="550" swimtime="00:12:19.46" />
                    <SPLIT distance="600" swimtime="00:13:29.71" />
                    <SPLIT distance="650" swimtime="00:14:38.80" />
                    <SPLIT distance="700" swimtime="00:15:47.42" />
                    <SPLIT distance="750" swimtime="00:16:56.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="118" swimtime="00:00:48.30" resultid="7566" heatid="10682" lane="8" entrytime="00:00:46.98" />
                <RESULT eventid="1226" points="137" swimtime="00:00:52.44" resultid="7567" heatid="10735" lane="4" entrytime="00:00:49.60" />
                <RESULT eventid="1287" points="100" swimtime="00:01:51.83" resultid="7568" heatid="10766" lane="8" entrytime="00:01:47.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="124" swimtime="00:01:56.48" resultid="7569" heatid="10840" lane="0" entrytime="00:01:58.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="93" swimtime="00:04:08.78" resultid="7570" heatid="10851" lane="5" entrytime="00:04:02.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.39" />
                    <SPLIT distance="100" swimtime="00:02:00.80" />
                    <SPLIT distance="150" swimtime="00:03:07.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="112" swimtime="00:04:16.65" resultid="7571" heatid="10894" lane="3" entrytime="00:04:08.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.06" />
                    <SPLIT distance="100" swimtime="00:02:06.27" />
                    <SPLIT distance="150" swimtime="00:03:14.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="90" swimtime="00:08:46.35" resultid="7572" heatid="10931" lane="7" entrytime="00:08:27.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.51" />
                    <SPLIT distance="100" swimtime="00:02:01.25" />
                    <SPLIT distance="150" swimtime="00:03:09.28" />
                    <SPLIT distance="200" swimtime="00:04:18.60" />
                    <SPLIT distance="250" swimtime="00:05:26.94" />
                    <SPLIT distance="300" swimtime="00:06:34.88" />
                    <SPLIT distance="350" swimtime="00:07:43.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-09-15" firstname="Adam" gender="M" lastname="Szmit" nation="POL" athleteid="5073">
              <RESULTS>
                <RESULT eventid="1128" points="224" swimtime="00:23:53.82" resultid="7605" heatid="10675" lane="3" entrytime="00:26:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                    <SPLIT distance="100" swimtime="00:01:25.19" />
                    <SPLIT distance="150" swimtime="00:02:12.01" />
                    <SPLIT distance="200" swimtime="00:02:59.66" />
                    <SPLIT distance="250" swimtime="00:03:46.69" />
                    <SPLIT distance="300" swimtime="00:04:34.89" />
                    <SPLIT distance="350" swimtime="00:05:21.86" />
                    <SPLIT distance="400" swimtime="00:06:09.28" />
                    <SPLIT distance="450" swimtime="00:06:57.22" />
                    <SPLIT distance="500" swimtime="00:07:46.03" />
                    <SPLIT distance="550" swimtime="00:08:34.40" />
                    <SPLIT distance="600" swimtime="00:09:22.75" />
                    <SPLIT distance="650" swimtime="00:10:11.43" />
                    <SPLIT distance="700" swimtime="00:10:59.76" />
                    <SPLIT distance="750" swimtime="00:11:42.08" />
                    <SPLIT distance="850" swimtime="00:13:21.74" />
                    <SPLIT distance="900" swimtime="00:14:13.81" />
                    <SPLIT distance="950" swimtime="00:15:02.52" />
                    <SPLIT distance="1000" swimtime="00:15:51.27" />
                    <SPLIT distance="1050" swimtime="00:16:39.24" />
                    <SPLIT distance="1100" swimtime="00:17:28.17" />
                    <SPLIT distance="1150" swimtime="00:18:17.10" />
                    <SPLIT distance="1200" swimtime="00:19:05.84" />
                    <SPLIT distance="1250" swimtime="00:19:55.46" />
                    <SPLIT distance="1300" swimtime="00:20:43.39" />
                    <SPLIT distance="1350" swimtime="00:21:27.08" />
                    <SPLIT distance="1400" swimtime="00:22:20.77" />
                    <SPLIT distance="1450" swimtime="00:23:03.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="240" swimtime="00:00:33.63" resultid="7606" heatid="10694" lane="0" entrytime="00:00:37.00" />
                <RESULT eventid="1302" points="244" swimtime="00:01:14.99" resultid="7607" heatid="10776" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="221" swimtime="00:02:48.70" resultid="7608" heatid="10859" lane="2" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:19.89" />
                    <SPLIT distance="150" swimtime="00:02:04.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="236" swimtime="00:05:55.82" resultid="7609" heatid="10939" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                    <SPLIT distance="100" swimtime="00:01:22.27" />
                    <SPLIT distance="150" swimtime="00:02:07.71" />
                    <SPLIT distance="200" swimtime="00:02:53.71" />
                    <SPLIT distance="250" swimtime="00:03:39.49" />
                    <SPLIT distance="300" swimtime="00:04:25.04" />
                    <SPLIT distance="350" swimtime="00:05:11.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-01" firstname="Gzegorz" gender="M" lastname="Mówiński" nation="POL" athleteid="5093">
              <RESULTS>
                <RESULT eventid="1128" points="219" swimtime="00:24:03.02" resultid="7622" heatid="10676" lane="0" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:27.75" />
                    <SPLIT distance="150" swimtime="00:02:15.21" />
                    <SPLIT distance="200" swimtime="00:03:03.30" />
                    <SPLIT distance="250" swimtime="00:03:50.67" />
                    <SPLIT distance="300" swimtime="00:04:39.13" />
                    <SPLIT distance="350" swimtime="00:05:27.14" />
                    <SPLIT distance="400" swimtime="00:06:15.76" />
                    <SPLIT distance="450" swimtime="00:07:04.58" />
                    <SPLIT distance="500" swimtime="00:07:53.03" />
                    <SPLIT distance="550" swimtime="00:08:41.69" />
                    <SPLIT distance="600" swimtime="00:09:30.15" />
                    <SPLIT distance="650" swimtime="00:10:18.53" />
                    <SPLIT distance="700" swimtime="00:11:07.74" />
                    <SPLIT distance="750" swimtime="00:11:56.20" />
                    <SPLIT distance="800" swimtime="00:12:45.10" />
                    <SPLIT distance="850" swimtime="00:13:33.29" />
                    <SPLIT distance="900" swimtime="00:14:22.53" />
                    <SPLIT distance="950" swimtime="00:15:10.90" />
                    <SPLIT distance="1000" swimtime="00:15:59.73" />
                    <SPLIT distance="1050" swimtime="00:16:48.03" />
                    <SPLIT distance="1100" swimtime="00:17:36.62" />
                    <SPLIT distance="1150" swimtime="00:18:25.11" />
                    <SPLIT distance="1200" swimtime="00:19:14.81" />
                    <SPLIT distance="1250" swimtime="00:20:03.18" />
                    <SPLIT distance="1300" swimtime="00:20:52.45" />
                    <SPLIT distance="1350" swimtime="00:21:41.72" />
                    <SPLIT distance="1400" swimtime="00:22:30.99" />
                    <SPLIT distance="1450" swimtime="00:23:18.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="184" swimtime="00:03:15.75" resultid="7623" heatid="10793" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:31.97" />
                    <SPLIT distance="150" swimtime="00:02:24.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="195" swimtime="00:07:00.40" resultid="7624" heatid="10877" lane="5" entrytime="00:07:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                    <SPLIT distance="100" swimtime="00:01:33.87" />
                    <SPLIT distance="150" swimtime="00:02:33.99" />
                    <SPLIT distance="200" swimtime="00:03:32.14" />
                    <SPLIT distance="250" swimtime="00:04:31.10" />
                    <SPLIT distance="300" swimtime="00:05:28.20" />
                    <SPLIT distance="350" swimtime="00:06:15.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="229" swimtime="00:05:59.19" resultid="7625" heatid="10939" lane="1" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                    <SPLIT distance="100" swimtime="00:01:25.45" />
                    <SPLIT distance="150" swimtime="00:02:12.13" />
                    <SPLIT distance="200" swimtime="00:02:59.24" />
                    <SPLIT distance="250" swimtime="00:03:45.86" />
                    <SPLIT distance="300" swimtime="00:04:32.41" />
                    <SPLIT distance="350" swimtime="00:05:17.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-25" firstname="Piotr" gender="M" lastname="Markowicz" nation="POL" athleteid="5045">
              <RESULTS>
                <RESULT eventid="1098" points="279" swimtime="00:11:31.21" resultid="7581" heatid="10672" lane="6" entrytime="00:10:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                    <SPLIT distance="100" swimtime="00:01:16.50" />
                    <SPLIT distance="150" swimtime="00:01:57.36" />
                    <SPLIT distance="200" swimtime="00:02:38.75" />
                    <SPLIT distance="250" swimtime="00:03:20.51" />
                    <SPLIT distance="300" swimtime="00:04:02.83" />
                    <SPLIT distance="350" swimtime="00:04:45.39" />
                    <SPLIT distance="400" swimtime="00:05:28.46" />
                    <SPLIT distance="450" swimtime="00:06:12.30" />
                    <SPLIT distance="500" swimtime="00:06:55.90" />
                    <SPLIT distance="550" swimtime="00:07:40.50" />
                    <SPLIT distance="600" swimtime="00:08:25.78" />
                    <SPLIT distance="650" swimtime="00:09:12.21" />
                    <SPLIT distance="700" swimtime="00:09:59.30" />
                    <SPLIT distance="750" swimtime="00:10:46.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="307" swimtime="00:00:30.99" resultid="7582" heatid="10701" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1190" points="276" swimtime="00:02:55.05" resultid="7583" heatid="10725" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                    <SPLIT distance="150" swimtime="00:02:15.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="7584" heatid="10747" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="337" swimtime="00:01:07.35" resultid="7585" heatid="10779" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="328" swimtime="00:00:32.52" resultid="7586" heatid="10832" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1482" points="311" swimtime="00:02:30.43" resultid="7587" heatid="10862" lane="9" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:13.37" />
                    <SPLIT distance="150" swimtime="00:01:51.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="290" swimtime="00:01:15.26" resultid="7588" heatid="10889" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="309" swimtime="00:05:25.41" resultid="7589" heatid="10942" lane="8" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:16.46" />
                    <SPLIT distance="150" swimtime="00:01:57.16" />
                    <SPLIT distance="200" swimtime="00:02:38.63" />
                    <SPLIT distance="250" swimtime="00:03:20.58" />
                    <SPLIT distance="300" swimtime="00:04:02.47" />
                    <SPLIT distance="350" swimtime="00:04:44.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-04-01" firstname="Piotr" gender="M" lastname="Konopacki" nation="POL" athleteid="5111">
              <RESULTS>
                <RESULT eventid="1098" points="345" swimtime="00:10:44.16" resultid="7637" heatid="10672" lane="5" entrytime="00:10:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:16.30" />
                    <SPLIT distance="150" swimtime="00:01:56.86" />
                    <SPLIT distance="200" swimtime="00:02:37.31" />
                    <SPLIT distance="250" swimtime="00:03:18.55" />
                    <SPLIT distance="300" swimtime="00:04:00.13" />
                    <SPLIT distance="350" swimtime="00:04:41.47" />
                    <SPLIT distance="400" swimtime="00:05:23.41" />
                    <SPLIT distance="450" swimtime="00:06:04.14" />
                    <SPLIT distance="500" swimtime="00:06:44.92" />
                    <SPLIT distance="550" swimtime="00:07:25.33" />
                    <SPLIT distance="600" swimtime="00:08:05.53" />
                    <SPLIT distance="650" swimtime="00:08:45.23" />
                    <SPLIT distance="700" swimtime="00:09:25.62" />
                    <SPLIT distance="750" swimtime="00:10:05.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="392" swimtime="00:00:28.56" resultid="7638" heatid="10703" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1302" points="385" swimtime="00:01:04.44" resultid="7639" heatid="10782" lane="1" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="357" swimtime="00:02:23.74" resultid="7640" heatid="10863" lane="0" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:08.68" />
                    <SPLIT distance="150" swimtime="00:01:46.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="377" swimtime="00:05:04.39" resultid="7641" heatid="10943" lane="8" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:11.94" />
                    <SPLIT distance="150" swimtime="00:01:51.55" />
                    <SPLIT distance="200" swimtime="00:02:30.86" />
                    <SPLIT distance="250" swimtime="00:03:10.75" />
                    <SPLIT distance="300" swimtime="00:03:50.07" />
                    <SPLIT distance="350" swimtime="00:04:29.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-25" firstname="Adam" gender="M" lastname="Matusiak vel Matuszewski" nation="POL" athleteid="5148">
              <RESULTS>
                <RESULT eventid="1128" points="161" swimtime="00:26:38.40" resultid="7668" heatid="10676" lane="7" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                    <SPLIT distance="100" swimtime="00:01:34.42" />
                    <SPLIT distance="150" swimtime="00:02:27.63" />
                    <SPLIT distance="200" swimtime="00:03:20.60" />
                    <SPLIT distance="250" swimtime="00:04:15.11" />
                    <SPLIT distance="300" swimtime="00:05:09.31" />
                    <SPLIT distance="350" swimtime="00:06:03.63" />
                    <SPLIT distance="400" swimtime="00:06:57.50" />
                    <SPLIT distance="450" swimtime="00:07:51.63" />
                    <SPLIT distance="500" swimtime="00:08:45.46" />
                    <SPLIT distance="550" swimtime="00:09:40.11" />
                    <SPLIT distance="600" swimtime="00:10:34.18" />
                    <SPLIT distance="650" swimtime="00:11:28.78" />
                    <SPLIT distance="700" swimtime="00:12:22.30" />
                    <SPLIT distance="750" swimtime="00:13:16.05" />
                    <SPLIT distance="800" swimtime="00:14:09.87" />
                    <SPLIT distance="850" swimtime="00:15:04.91" />
                    <SPLIT distance="900" swimtime="00:15:58.93" />
                    <SPLIT distance="950" swimtime="00:16:54.20" />
                    <SPLIT distance="1000" swimtime="00:17:47.73" />
                    <SPLIT distance="1050" swimtime="00:18:42.60" />
                    <SPLIT distance="1100" swimtime="00:19:36.43" />
                    <SPLIT distance="1150" swimtime="00:20:31.46" />
                    <SPLIT distance="1200" swimtime="00:21:25.02" />
                    <SPLIT distance="1250" swimtime="00:22:19.94" />
                    <SPLIT distance="1350" swimtime="00:22:36.29" />
                    <SPLIT distance="1400" swimtime="00:23:14.31" />
                    <SPLIT distance="1450" swimtime="00:23:29.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="207" swimtime="00:00:35.34" resultid="7669" heatid="10695" lane="0" entrytime="00:00:35.12" />
                <RESULT eventid="1242" points="136" swimtime="00:00:46.68" resultid="7670" heatid="10740" lane="6" />
                <RESULT eventid="1302" points="195" swimtime="00:01:20.89" resultid="7671" heatid="10776" lane="1" entrytime="00:01:19.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="139" swimtime="00:00:43.28" resultid="7672" heatid="10827" lane="4" entrytime="00:00:42.89" />
                <RESULT eventid="1482" points="190" swimtime="00:02:57.40" resultid="7673" heatid="10859" lane="7" entrytime="00:02:54.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:25.80" />
                    <SPLIT distance="150" swimtime="00:02:12.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="7674" heatid="10900" lane="7" entrytime="00:03:40.21" />
                <RESULT eventid="1695" points="176" swimtime="00:06:32.18" resultid="7675" heatid="10938" lane="0" entrytime="00:06:30.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                    <SPLIT distance="100" swimtime="00:01:34.12" />
                    <SPLIT distance="150" swimtime="00:02:25.79" />
                    <SPLIT distance="200" swimtime="00:03:17.21" />
                    <SPLIT distance="250" swimtime="00:04:08.75" />
                    <SPLIT distance="300" swimtime="00:04:59.98" />
                    <SPLIT distance="350" swimtime="00:05:49.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-16" firstname="Paweł" gender="M" lastname="Szczuka" nation="POL" athleteid="5068">
              <RESULTS>
                <RESULT eventid="1190" points="444" swimtime="00:02:29.33" resultid="7601" heatid="10729" lane="6" entrytime="00:02:28.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                    <SPLIT distance="150" swimtime="00:01:55.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="430" swimtime="00:00:31.85" resultid="7602" heatid="10750" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1452" points="363" swimtime="00:01:12.66" resultid="7603" heatid="10848" lane="7" entrytime="00:01:15.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="444" swimtime="00:05:19.54" resultid="7604" heatid="10880" lane="5" entrytime="00:05:29.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="150" swimtime="00:01:51.89" />
                    <SPLIT distance="200" swimtime="00:02:35.22" />
                    <SPLIT distance="250" swimtime="00:03:21.57" />
                    <SPLIT distance="300" swimtime="00:04:07.44" />
                    <SPLIT distance="350" swimtime="00:04:43.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="5117">
              <RESULTS>
                <RESULT eventid="1098" points="460" swimtime="00:09:45.58" resultid="7642" heatid="10673" lane="7" entrytime="00:09:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="150" swimtime="00:01:45.87" />
                    <SPLIT distance="200" swimtime="00:02:22.88" />
                    <SPLIT distance="250" swimtime="00:02:59.93" />
                    <SPLIT distance="300" swimtime="00:03:37.02" />
                    <SPLIT distance="350" swimtime="00:04:14.24" />
                    <SPLIT distance="400" swimtime="00:04:51.31" />
                    <SPLIT distance="450" swimtime="00:05:28.17" />
                    <SPLIT distance="500" swimtime="00:06:04.89" />
                    <SPLIT distance="550" swimtime="00:06:42.00" />
                    <SPLIT distance="600" swimtime="00:07:18.94" />
                    <SPLIT distance="650" swimtime="00:07:55.84" />
                    <SPLIT distance="700" swimtime="00:08:32.64" />
                    <SPLIT distance="750" swimtime="00:09:09.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="474" swimtime="00:00:26.80" resultid="7643" heatid="10706" lane="3" entrytime="00:00:27.50" />
                <RESULT eventid="1190" points="418" swimtime="00:02:32.40" resultid="7644" heatid="10729" lane="1" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="100" swimtime="00:01:13.90" />
                    <SPLIT distance="150" swimtime="00:01:58.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="527" swimtime="00:00:58.07" resultid="7645" heatid="10786" lane="2" entrytime="00:00:58.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="484" swimtime="00:02:09.85" resultid="7646" heatid="10866" lane="9" entrytime="00:02:09.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                    <SPLIT distance="150" swimtime="00:01:38.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="391" swimtime="00:05:33.27" resultid="7647" heatid="10880" lane="6" entrytime="00:05:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:58.79" />
                    <SPLIT distance="200" swimtime="00:02:43.74" />
                    <SPLIT distance="250" swimtime="00:03:32.87" />
                    <SPLIT distance="300" swimtime="00:04:19.28" />
                    <SPLIT distance="350" swimtime="00:04:56.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="7648" heatid="10890" lane="4" entrytime="00:01:05.60" />
                <RESULT eventid="1695" points="492" swimtime="00:04:38.74" resultid="7649" heatid="10944" lane="5" entrytime="00:04:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="100" swimtime="00:01:07.14" />
                    <SPLIT distance="150" swimtime="00:01:42.32" />
                    <SPLIT distance="200" swimtime="00:02:18.33" />
                    <SPLIT distance="250" swimtime="00:02:53.95" />
                    <SPLIT distance="300" swimtime="00:03:29.66" />
                    <SPLIT distance="350" swimtime="00:04:05.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-29" firstname="Jakub" gender="M" lastname="Stępień" nation="POL" athleteid="5079">
              <RESULTS>
                <RESULT eventid="1128" points="219" swimtime="00:24:03.74" resultid="7610" heatid="10678" lane="1" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:01:23.63" />
                    <SPLIT distance="150" swimtime="00:02:09.83" />
                    <SPLIT distance="200" swimtime="00:02:57.11" />
                    <SPLIT distance="250" swimtime="00:03:46.21" />
                    <SPLIT distance="300" swimtime="00:04:35.96" />
                    <SPLIT distance="350" swimtime="00:05:24.88" />
                    <SPLIT distance="400" swimtime="00:06:14.14" />
                    <SPLIT distance="450" swimtime="00:07:03.14" />
                    <SPLIT distance="500" swimtime="00:07:52.52" />
                    <SPLIT distance="550" swimtime="00:08:41.50" />
                    <SPLIT distance="600" swimtime="00:09:31.13" />
                    <SPLIT distance="650" swimtime="00:10:20.90" />
                    <SPLIT distance="700" swimtime="00:11:10.47" />
                    <SPLIT distance="750" swimtime="00:11:59.88" />
                    <SPLIT distance="800" swimtime="00:12:49.72" />
                    <SPLIT distance="850" swimtime="00:13:39.53" />
                    <SPLIT distance="900" swimtime="00:14:29.42" />
                    <SPLIT distance="950" swimtime="00:15:18.52" />
                    <SPLIT distance="1000" swimtime="00:16:07.78" />
                    <SPLIT distance="1050" swimtime="00:16:56.47" />
                    <SPLIT distance="1100" swimtime="00:17:44.70" />
                    <SPLIT distance="1150" swimtime="00:18:32.85" />
                    <SPLIT distance="1200" swimtime="00:19:21.03" />
                    <SPLIT distance="1250" swimtime="00:20:09.14" />
                    <SPLIT distance="1300" swimtime="00:20:57.20" />
                    <SPLIT distance="1350" swimtime="00:21:44.28" />
                    <SPLIT distance="1400" swimtime="00:22:31.73" />
                    <SPLIT distance="1450" swimtime="00:23:19.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="338" swimtime="00:00:30.00" resultid="7611" heatid="10703" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="7612" heatid="10781" lane="2" entrytime="00:01:05.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="7613" heatid="10831" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1482" points="308" swimtime="00:02:31.00" resultid="7614" heatid="10862" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:10.09" />
                    <SPLIT distance="150" swimtime="00:01:51.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="5085">
              <RESULTS>
                <RESULT eventid="1098" points="346" swimtime="00:10:43.93" resultid="7615" heatid="10668" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:16.53" />
                    <SPLIT distance="150" swimtime="00:01:57.09" />
                    <SPLIT distance="200" swimtime="00:02:37.71" />
                    <SPLIT distance="250" swimtime="00:03:18.69" />
                    <SPLIT distance="300" swimtime="00:03:59.58" />
                    <SPLIT distance="350" swimtime="00:04:40.67" />
                    <SPLIT distance="400" swimtime="00:05:21.40" />
                    <SPLIT distance="450" swimtime="00:06:02.39" />
                    <SPLIT distance="500" swimtime="00:06:43.00" />
                    <SPLIT distance="550" swimtime="00:07:23.94" />
                    <SPLIT distance="600" swimtime="00:08:04.70" />
                    <SPLIT distance="650" swimtime="00:08:45.68" />
                    <SPLIT distance="700" swimtime="00:09:26.54" />
                    <SPLIT distance="750" swimtime="00:10:06.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="7616" heatid="10724" lane="7" entrytime="00:02:55.00" />
                <RESULT eventid="1332" points="234" swimtime="00:03:00.73" resultid="7617" heatid="10795" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:26.83" />
                    <SPLIT distance="150" swimtime="00:02:14.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="337" swimtime="00:00:32.22" resultid="7618" heatid="10829" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1546" status="DNS" swimtime="00:00:00.00" resultid="7619" heatid="10879" lane="8" entrytime="00:06:15.00" />
                <RESULT eventid="1578" points="324" swimtime="00:01:12.47" resultid="7620" heatid="10888" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="338" swimtime="00:05:15.72" resultid="7621" heatid="10940" lane="5" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:18.55" />
                    <SPLIT distance="150" swimtime="00:01:59.00" />
                    <SPLIT distance="200" swimtime="00:02:39.41" />
                    <SPLIT distance="250" swimtime="00:03:19.79" />
                    <SPLIT distance="300" swimtime="00:03:59.85" />
                    <SPLIT distance="350" swimtime="00:04:39.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-02-09" firstname="Aleksandra" gender="F" lastname="Milewska" nation="POL" athleteid="5142">
              <RESULTS>
                <RESULT eventid="1175" points="347" swimtime="00:02:59.39" resultid="7663" heatid="10716" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:01:25.13" />
                    <SPLIT distance="150" swimtime="00:02:16.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" status="DNS" swimtime="00:00:00.00" resultid="7664" heatid="10737" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1287" points="390" swimtime="00:01:11.21" resultid="7665" heatid="10769" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="369" swimtime="00:00:34.03" resultid="7666" heatid="10823" lane="2" entrytime="00:00:34.50" />
                <RESULT eventid="1467" points="342" swimtime="00:02:41.54" resultid="7667" heatid="10854" lane="3" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                    <SPLIT distance="150" swimtime="00:01:59.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-13" firstname="Michał" gender="M" lastname="Kieres" nation="POL" athleteid="5098">
              <RESULTS>
                <RESULT eventid="1190" points="305" swimtime="00:02:49.31" resultid="7626" heatid="10725" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:21.14" />
                    <SPLIT distance="150" swimtime="00:02:09.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="341" swimtime="00:03:01.67" resultid="7627" heatid="10763" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:23.96" />
                    <SPLIT distance="150" swimtime="00:02:12.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="285" swimtime="00:02:49.42" resultid="7628" heatid="10795" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:02:02.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="306" swimtime="00:06:01.50" resultid="7630" heatid="10880" lane="4" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:02:06.98" />
                    <SPLIT distance="200" swimtime="00:02:58.02" />
                    <SPLIT distance="250" swimtime="00:03:47.74" />
                    <SPLIT distance="300" swimtime="00:04:38.27" />
                    <SPLIT distance="350" swimtime="00:05:20.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="313" swimtime="00:01:13.32" resultid="7631" heatid="10890" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="374" swimtime="00:00:36.64" resultid="7632" heatid="10921" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1392" points="345" swimtime="00:01:21.39" resultid="10612" heatid="10817" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-10-03" firstname="Bartosz" gender="M" lastname="Wolak" nation="POL" athleteid="5062">
              <RESULTS>
                <RESULT eventid="1160" points="482" swimtime="00:00:26.66" resultid="7596" heatid="10707" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1302" points="455" swimtime="00:01:00.96" resultid="7597" heatid="10784" lane="2" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="438" swimtime="00:00:29.53" resultid="7598" heatid="10835" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="1482" points="361" swimtime="00:02:23.23" resultid="7599" heatid="10864" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:07.81" />
                    <SPLIT distance="150" swimtime="00:01:45.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="408" swimtime="00:01:07.16" resultid="7600" heatid="10890" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-06-26" firstname="Monika" gender="F" lastname="Piwońska" nation="POL" athleteid="5157">
              <RESULTS>
                <RESULT eventid="1113" points="299" swimtime="00:23:02.68" resultid="7676" heatid="10674" lane="6" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:21.84" />
                    <SPLIT distance="150" swimtime="00:02:07.08" />
                    <SPLIT distance="200" swimtime="00:02:52.69" />
                    <SPLIT distance="250" swimtime="00:03:38.11" />
                    <SPLIT distance="300" swimtime="00:04:23.75" />
                    <SPLIT distance="350" swimtime="00:05:09.76" />
                    <SPLIT distance="400" swimtime="00:05:55.98" />
                    <SPLIT distance="450" swimtime="00:06:41.87" />
                    <SPLIT distance="500" swimtime="00:07:28.14" />
                    <SPLIT distance="550" swimtime="00:08:14.94" />
                    <SPLIT distance="600" swimtime="00:09:01.96" />
                    <SPLIT distance="650" swimtime="00:09:48.81" />
                    <SPLIT distance="700" swimtime="00:10:35.83" />
                    <SPLIT distance="750" swimtime="00:11:22.53" />
                    <SPLIT distance="800" swimtime="00:12:09.36" />
                    <SPLIT distance="850" swimtime="00:12:56.37" />
                    <SPLIT distance="900" swimtime="00:13:43.28" />
                    <SPLIT distance="950" swimtime="00:14:30.49" />
                    <SPLIT distance="1000" swimtime="00:15:17.52" />
                    <SPLIT distance="1050" swimtime="00:16:04.30" />
                    <SPLIT distance="1100" swimtime="00:16:51.18" />
                    <SPLIT distance="1150" swimtime="00:17:38.56" />
                    <SPLIT distance="1200" swimtime="00:18:25.91" />
                    <SPLIT distance="1250" swimtime="00:19:13.02" />
                    <SPLIT distance="1300" swimtime="00:19:59.24" />
                    <SPLIT distance="1350" swimtime="00:20:44.77" />
                    <SPLIT distance="1400" swimtime="00:21:31.38" />
                    <SPLIT distance="1450" swimtime="00:22:17.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="414" swimtime="00:02:49.21" resultid="7677" heatid="10717" lane="6" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:18.95" />
                    <SPLIT distance="150" swimtime="00:02:09.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1317" points="287" swimtime="00:03:04.56" resultid="7678" heatid="10790" lane="4" entrytime="00:02:58.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="100" swimtime="00:01:27.54" />
                    <SPLIT distance="150" swimtime="00:02:17.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="428" swimtime="00:00:32.41" resultid="7679" heatid="10824" lane="0" entrytime="00:00:33.23" />
                <RESULT eventid="1525" points="367" swimtime="00:06:11.78" resultid="7680" heatid="10875" lane="8" entrytime="00:06:01.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:22.34" />
                    <SPLIT distance="150" swimtime="00:02:13.69" />
                    <SPLIT distance="200" swimtime="00:03:01.35" />
                    <SPLIT distance="250" swimtime="00:03:52.73" />
                    <SPLIT distance="300" swimtime="00:04:42.95" />
                    <SPLIT distance="350" swimtime="00:05:27.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-14" firstname="Wojciech" gender="M" lastname="Kłujszo" nation="POL" athleteid="5126">
              <RESULTS>
                <RESULT eventid="1160" points="292" swimtime="00:00:31.51" resultid="7650" heatid="10698" lane="6" entrytime="00:00:31.70" />
                <RESULT eventid="1638" points="272" swimtime="00:00:40.73" resultid="7651" heatid="10917" lane="6" entrytime="00:00:40.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-26" firstname="Joanna" gender="F" lastname="Drzewicka" nation="POL" athleteid="5129">
              <RESULTS>
                <RESULT eventid="1059" points="176" swimtime="00:14:24.92" resultid="7652" heatid="10665" lane="3" />
                <RESULT eventid="1144" points="273" swimtime="00:00:36.55" resultid="7653" heatid="10683" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="7654" heatid="10714" lane="5" entrytime="00:03:30.00" />
                <RESULT eventid="1226" points="308" swimtime="00:00:40.04" resultid="7655" heatid="10737" lane="6" entrytime="00:00:40.30" />
                <RESULT eventid="1287" points="224" swimtime="00:01:25.72" resultid="7656" heatid="10767" lane="3" entrytime="00:01:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="268" swimtime="00:01:30.11" resultid="7657" heatid="10841" lane="9" entrytime="00:01:30.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="230" swimtime="00:03:22.24" resultid="7658" heatid="10895" lane="6" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.94" />
                    <SPLIT distance="100" swimtime="00:01:40.41" />
                    <SPLIT distance="150" swimtime="00:02:32.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="Kucharska" nation="POL" athleteid="5137">
              <RESULTS>
                <RESULT eventid="1144" points="359" swimtime="00:00:33.37" resultid="7659" heatid="10685" lane="4" entrytime="00:00:33.80" />
                <RESULT eventid="1226" points="307" swimtime="00:00:40.08" resultid="7660" heatid="10737" lane="2" entrytime="00:00:40.50" />
                <RESULT eventid="1287" points="326" swimtime="00:01:15.59" resultid="7661" heatid="10769" lane="0" entrytime="00:01:16.50" />
                <RESULT eventid="1593" points="257" swimtime="00:03:14.92" resultid="7662" heatid="10896" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                    <SPLIT distance="100" swimtime="00:01:34.86" />
                    <SPLIT distance="150" swimtime="00:02:26.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-09" firstname="Marek" gender="M" lastname="Koźlikowski" nation="POL" athleteid="5038">
              <RESULTS>
                <RESULT eventid="1128" status="DNS" swimtime="00:00:00.00" resultid="7575" heatid="10676" lane="1" entrytime="00:25:00.00" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="7576" heatid="10721" lane="3" entrytime="00:03:25.23" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="7577" heatid="10759" lane="2" entrytime="00:03:30.22" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="7578" heatid="10828" lane="0" entrytime="00:00:40.23" />
                <RESULT eventid="1546" status="DNS" swimtime="00:00:00.00" resultid="7579" heatid="10877" lane="4" entrytime="00:07:00.23" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="7580" heatid="10939" lane="5" entrytime="00:06:00.25" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="321" swimtime="00:02:16.44" resultid="7683" heatid="10801" lane="8" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="100" swimtime="00:01:13.22" />
                    <SPLIT distance="150" swimtime="00:01:45.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5085" number="1" />
                    <RELAYPOSITION athleteid="5098" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5045" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5106" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" points="320" swimtime="00:02:03.94" resultid="7686" heatid="10871" lane="2" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:02.39" />
                    <SPLIT distance="150" swimtime="00:01:32.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5106" number="1" />
                    <RELAYPOSITION athleteid="5045" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5079" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5085" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1368" points="483" swimtime="00:01:59.00" resultid="7681" heatid="10802" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                    <SPLIT distance="150" swimtime="00:01:32.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5111" number="1" />
                    <RELAYPOSITION athleteid="5068" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5055" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5117" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" points="512" swimtime="00:01:46.01" resultid="7682" heatid="10872" lane="6" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                    <SPLIT distance="100" swimtime="00:00:54.70" />
                    <SPLIT distance="150" swimtime="00:01:21.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5068" number="1" />
                    <RELAYPOSITION athleteid="5117" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5111" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5055" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1518" status="DNS" swimtime="00:00:00.00" resultid="7687" heatid="10870" lane="3" entrytime="00:02:06.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5098" number="1" />
                    <RELAYPOSITION athleteid="5038" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5093" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5126" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1368" status="DNS" swimtime="00:00:00.00" resultid="7684" heatid="10800" lane="5" entrytime="00:02:29.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5148" number="1" />
                    <RELAYPOSITION athleteid="5093" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5038" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5073" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1368" status="DNS" swimtime="00:00:00.00" resultid="7689" heatid="10802" lane="6" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5111" number="1" />
                    <RELAYPOSITION athleteid="5068" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5055" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5117" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:01:59.54" resultid="7685" heatid="10733" lane="9" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.14" />
                    <SPLIT distance="100" swimtime="00:01:00.62" />
                    <SPLIT distance="150" swimtime="00:01:33.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5055" number="1" />
                    <RELAYPOSITION athleteid="5129" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5137" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5068" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:14.50" resultid="7688" heatid="10929" lane="9" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:15.01" />
                    <SPLIT distance="150" swimtime="00:01:41.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5129" number="1" />
                    <RELAYPOSITION athleteid="5117" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5055" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5137" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AQGDY" nation="POL" region="07" clubid="10611" name="AquaStars Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1978-01-01" firstname="Mariusz" gender="M" lastname="Golon" nation="POL" athleteid="9768">
              <RESULTS>
                <RESULT eventid="1272" points="247" swimtime="00:03:22.23" resultid="10560" heatid="10760" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:37.12" />
                    <SPLIT distance="150" swimtime="00:02:32.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="10561" heatid="10810" lane="5" entrytime="00:01:50.00" />
                <RESULT eventid="1422" points="459" swimtime="00:00:29.07" resultid="10562" heatid="10832" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1638" points="434" swimtime="00:00:34.87" resultid="10563" heatid="10918" lane="9" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZS UW" nation="POL" region="MAZ" clubid="3054" name="AZS  Klub Uczelniany Uniwersytetu Warszawskiego" shortname="AZS  Klub Uczelniany Uniwersyt">
          <CONTACT city="Warszawa" email="mbaranowski@biogeo.uw.edu.pl, azs@uw.edu.pl," internet="www.kuazsuw.pl" name="Baranowski Marek" phone="602445201" state="MAZ" street="Krakowskie Przedmieście" zip="00-325" />
          <ATHLETES>
            <ATHLETE birthdate="1991-01-15" firstname="Marek" gender="M" lastname="Baranowski" nation="POL" athleteid="3055">
              <RESULTS>
                <RESULT eventid="1302" points="539" swimtime="00:00:57.63" resultid="8437" heatid="10786" lane="3" entrytime="00:00:58.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="454" swimtime="00:02:12.65" resultid="8438" heatid="10866" lane="4" entrytime="00:02:14.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                    <SPLIT distance="100" swimtime="00:01:01.43" />
                    <SPLIT distance="150" swimtime="00:01:36.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" region="11" clubid="3156" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501 370 222" state="ŚLASK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1931-04-27" firstname="Jan" gender="M" lastname="Ślężyński" nation="POL" license="100611700315" athleteid="3157">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Mężczyzn  w  kat M 85-89  lat" eventid="1128" points="34" swimtime="00:44:33.69" resultid="3158" heatid="10675" lane="0" entrytime="00:47:50.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.08" />
                    <SPLIT distance="100" swimtime="00:02:36.66" />
                    <SPLIT distance="150" swimtime="00:04:01.27" />
                    <SPLIT distance="200" swimtime="00:05:30.34" />
                    <SPLIT distance="250" swimtime="00:06:57.61" />
                    <SPLIT distance="300" swimtime="00:08:25.56" />
                    <SPLIT distance="350" swimtime="00:09:54.52" />
                    <SPLIT distance="400" swimtime="00:11:24.30" />
                    <SPLIT distance="450" swimtime="00:12:51.71" />
                    <SPLIT distance="500" swimtime="00:14:22.82" />
                    <SPLIT distance="550" swimtime="00:15:52.54" />
                    <SPLIT distance="600" swimtime="00:17:24.21" />
                    <SPLIT distance="650" swimtime="00:18:54.06" />
                    <SPLIT distance="700" swimtime="00:20:24.48" />
                    <SPLIT distance="750" swimtime="00:21:55.28" />
                    <SPLIT distance="800" swimtime="00:23:27.43" />
                    <SPLIT distance="850" swimtime="00:24:57.65" />
                    <SPLIT distance="900" swimtime="00:26:29.06" />
                    <SPLIT distance="950" swimtime="00:27:59.69" />
                    <SPLIT distance="1000" swimtime="00:29:31.12" />
                    <SPLIT distance="1050" swimtime="00:31:02.41" />
                    <SPLIT distance="1100" swimtime="00:32:32.70" />
                    <SPLIT distance="1150" swimtime="00:34:02.61" />
                    <SPLIT distance="1200" swimtime="00:35:33.50" />
                    <SPLIT distance="1250" swimtime="00:37:04.73" />
                    <SPLIT distance="1300" swimtime="00:38:36.57" />
                    <SPLIT distance="1350" swimtime="00:40:08.18" />
                    <SPLIT distance="1400" swimtime="00:41:38.86" />
                    <SPLIT distance="1450" swimtime="00:43:08.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="45" swimtime="00:00:58.48" resultid="3159" heatid="10689" lane="0" entrytime="00:01:06.34" />
                <RESULT eventid="1272" points="39" swimtime="00:06:14.21" resultid="3160" heatid="10757" lane="3" entrytime="00:05:58.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.74" />
                    <SPLIT distance="100" swimtime="00:03:02.87" />
                    <SPLIT distance="150" swimtime="00:04:42.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="29" swimtime="00:02:32.20" resultid="3161" heatid="10773" lane="7" entrytime="00:02:30.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="36" swimtime="00:02:52.70" resultid="3162" heatid="10809" lane="3" entrytime="00:02:49.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="33" swimtime="00:05:15.41" resultid="3163" heatid="10856" lane="5" entrytime="00:05:36.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.68" />
                    <SPLIT distance="100" swimtime="00:02:36.17" />
                    <SPLIT distance="150" swimtime="00:04:00.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="46" swimtime="00:01:13.73" resultid="3164" heatid="10913" lane="0" entrytime="00:01:10.23" />
                <RESULT eventid="1695" points="35" swimtime="00:11:09.60" resultid="3165" heatid="10936" lane="0" entrytime="00:11:34.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.26" />
                    <SPLIT distance="100" swimtime="00:02:39.83" />
                    <SPLIT distance="150" swimtime="00:04:07.02" />
                    <SPLIT distance="200" swimtime="00:05:34.97" />
                    <SPLIT distance="250" swimtime="00:06:59.61" />
                    <SPLIT distance="300" swimtime="00:08:26.28" />
                    <SPLIT distance="350" swimtime="00:09:51.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZRAC" nation="POL" region="SLA" clubid="2956" name="AZS PWSZ Raciborz">
          <CONTACT city="Racibórz" email="adip45@poczta.onet.pl" name="M Kunicki" state="ŚL" street="słowackiego 55" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1957-04-11" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="2957">
              <RESULTS>
                <RESULT eventid="1190" points="226" swimtime="00:03:07.11" resultid="7922" heatid="10722" lane="7" entrytime="00:03:10.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:27.28" />
                    <SPLIT distance="150" swimtime="00:02:22.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="241" swimtime="00:03:23.92" resultid="7923" heatid="10760" lane="6" entrytime="00:03:19.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                    <SPLIT distance="100" swimtime="00:01:38.54" />
                    <SPLIT distance="150" swimtime="00:02:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="174" swimtime="00:03:19.61" resultid="7924" heatid="10793" lane="6" entrytime="00:03:15.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.28" />
                    <SPLIT distance="100" swimtime="00:01:34.72" />
                    <SPLIT distance="150" swimtime="00:02:27.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="250" swimtime="00:01:30.65" resultid="7925" heatid="10814" lane="9" entrytime="00:01:29.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="221" swimtime="00:06:42.78" resultid="7926" heatid="10878" lane="3" entrytime="00:06:38.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                    <SPLIT distance="100" swimtime="00:01:37.61" />
                    <SPLIT distance="150" swimtime="00:02:29.49" />
                    <SPLIT distance="200" swimtime="00:03:21.13" />
                    <SPLIT distance="250" swimtime="00:04:18.02" />
                    <SPLIT distance="300" swimtime="00:05:13.39" />
                    <SPLIT distance="350" swimtime="00:05:59.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="175" swimtime="00:01:28.94" resultid="7927" heatid="10887" lane="2" entrytime="00:01:25.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="297" swimtime="00:00:39.56" resultid="7928" heatid="10919" lane="1" entrytime="00:00:39.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CMMAS" nation="POL" region="14" clubid="9543" name="AZS UJ CM Masters">
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Jacek" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="6200">
              <RESULTS>
                <RESULT eventid="1128" points="198" swimtime="00:24:53.67" resultid="9542" heatid="10676" lane="8" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.22" />
                    <SPLIT distance="100" swimtime="00:01:32.60" />
                    <SPLIT distance="150" swimtime="00:02:22.33" />
                    <SPLIT distance="200" swimtime="00:03:12.06" />
                    <SPLIT distance="250" swimtime="00:04:01.52" />
                    <SPLIT distance="300" swimtime="00:04:51.96" />
                    <SPLIT distance="350" swimtime="00:05:41.98" />
                    <SPLIT distance="400" swimtime="00:06:31.29" />
                    <SPLIT distance="450" swimtime="00:07:21.28" />
                    <SPLIT distance="500" swimtime="00:08:12.60" />
                    <SPLIT distance="550" swimtime="00:09:02.46" />
                    <SPLIT distance="600" swimtime="00:09:54.09" />
                    <SPLIT distance="650" swimtime="00:10:44.56" />
                    <SPLIT distance="700" swimtime="00:11:35.01" />
                    <SPLIT distance="750" swimtime="00:12:24.02" />
                    <SPLIT distance="800" swimtime="00:13:15.35" />
                    <SPLIT distance="850" swimtime="00:14:05.71" />
                    <SPLIT distance="900" swimtime="00:14:54.55" />
                    <SPLIT distance="950" swimtime="00:15:45.63" />
                    <SPLIT distance="1000" swimtime="00:16:35.82" />
                    <SPLIT distance="1050" swimtime="00:17:26.27" />
                    <SPLIT distance="1100" swimtime="00:18:16.47" />
                    <SPLIT distance="1150" swimtime="00:19:06.31" />
                    <SPLIT distance="1200" swimtime="00:19:57.71" />
                    <SPLIT distance="1250" swimtime="00:20:48.24" />
                    <SPLIT distance="1300" swimtime="00:21:38.36" />
                    <SPLIT distance="1350" swimtime="00:22:27.65" />
                    <SPLIT distance="1400" swimtime="00:23:18.26" />
                    <SPLIT distance="1450" swimtime="00:24:08.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BABIA" nation="POL" region="PDL" clubid="5596" name="Barracuda Białystok">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1953-01-01" firstname="Mirosław" gender="M" lastname="Gawryluk" nation="POL" athleteid="5597">
              <RESULTS>
                <RESULT eventid="1160" points="138" swimtime="00:00:40.40" resultid="7105" heatid="10690" lane="1" />
                <RESULT eventid="1302" points="110" swimtime="00:01:37.66" resultid="7106" heatid="10772" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1368" status="DNS" swimtime="00:00:00.00" resultid="7117" heatid="10800" lane="4" entrytime="00:02:24.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5597" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" status="DNS" swimtime="00:00:00.00" resultid="7118" heatid="10871" lane="0" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5597" number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="BLGRO" nation="BLR" clubid="6122" name="BLR GRODNO &quot; MKTeam&quot;">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1950-01-01" firstname="Nadzeya" gender="F" lastname="Kuzmina" nation="BLR" athleteid="6197">
              <RESULTS>
                <RESULT eventid="1144" points="163" swimtime="00:00:43.39" resultid="7481" heatid="10682" lane="6" entrytime="00:00:43.50" />
                <RESULT eventid="1623" points="128" swimtime="00:00:58.48" resultid="7482" heatid="10906" lane="8" entrytime="00:01:00.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Yury" gender="M" lastname="Komov" nation="BLR" athleteid="6192">
              <RESULTS>
                <RESULT eventid="1160" points="230" swimtime="00:00:34.09" resultid="7477" heatid="10694" lane="3" entrytime="00:00:35.20" />
                <RESULT eventid="1272" points="220" swimtime="00:03:30.29" resultid="7478" heatid="10759" lane="8" entrytime="00:03:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.04" />
                    <SPLIT distance="100" swimtime="00:01:38.17" />
                    <SPLIT distance="150" swimtime="00:02:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="249" swimtime="00:01:30.74" resultid="7479" heatid="10812" lane="2" entrytime="00:01:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="324" swimtime="00:00:38.45" resultid="7480" heatid="10917" lane="8" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ACWRO" nation="POL" region="DOL" clubid="9320" name="Fitness Academy Wrocław">
          <CONTACT city="Wrocław" name="Wolny Dariusz" phone="603630870" state="DOL" street="Rogowska 52a" zip="54-440" />
          <ATHLETES>
            <ATHLETE birthdate="1960-05-11" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="9350">
              <RESULTS>
                <RESULT eventid="1175" points="168" swimtime="00:03:48.43" resultid="9351" heatid="10714" lane="8" entrytime="00:03:47.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.58" />
                    <SPLIT distance="100" swimtime="00:01:56.80" />
                    <SPLIT distance="150" swimtime="00:02:58.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="217" swimtime="00:03:51.45" resultid="9352" heatid="10754" lane="2" entrytime="00:03:47.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.41" />
                    <SPLIT distance="100" swimtime="00:01:51.34" />
                    <SPLIT distance="150" swimtime="00:02:52.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="190" swimtime="00:01:30.40" resultid="9353" heatid="10767" lane="6" entrytime="00:01:26.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="233" swimtime="00:01:44.48" resultid="9354" heatid="10805" lane="2" entrytime="00:01:42.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="122" swimtime="00:00:49.19" resultid="9355" heatid="10821" lane="1" entrytime="00:00:47.59" />
                <RESULT eventid="1623" points="236" swimtime="00:00:47.69" resultid="9356" heatid="10908" lane="1" entrytime="00:00:45.77" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-13" firstname="Małgorzata" gender="F" lastname="Bołtuć" nation="POL" athleteid="9343">
              <RESULTS>
                <RESULT eventid="1113" points="217" swimtime="00:25:38.34" resultid="9344" heatid="10674" lane="7" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                    <SPLIT distance="100" swimtime="00:01:34.74" />
                    <SPLIT distance="150" swimtime="00:02:24.67" />
                    <SPLIT distance="200" swimtime="00:03:15.31" />
                    <SPLIT distance="250" swimtime="00:04:06.26" />
                    <SPLIT distance="300" swimtime="00:04:58.32" />
                    <SPLIT distance="350" swimtime="00:05:49.43" />
                    <SPLIT distance="400" swimtime="00:06:40.32" />
                    <SPLIT distance="450" swimtime="00:07:32.07" />
                    <SPLIT distance="500" swimtime="00:08:23.80" />
                    <SPLIT distance="550" swimtime="00:09:15.22" />
                    <SPLIT distance="600" swimtime="00:10:07.32" />
                    <SPLIT distance="650" swimtime="00:10:58.40" />
                    <SPLIT distance="700" swimtime="00:11:49.90" />
                    <SPLIT distance="750" swimtime="00:12:41.05" />
                    <SPLIT distance="800" swimtime="00:13:32.66" />
                    <SPLIT distance="850" swimtime="00:14:23.95" />
                    <SPLIT distance="900" swimtime="00:15:16.13" />
                    <SPLIT distance="950" swimtime="00:16:08.06" />
                    <SPLIT distance="1000" swimtime="00:17:00.87" />
                    <SPLIT distance="1050" swimtime="00:17:53.42" />
                    <SPLIT distance="1100" swimtime="00:18:45.16" />
                    <SPLIT distance="1150" swimtime="00:19:37.07" />
                    <SPLIT distance="1200" swimtime="00:20:29.29" />
                    <SPLIT distance="1250" swimtime="00:21:21.53" />
                    <SPLIT distance="1300" swimtime="00:22:13.64" />
                    <SPLIT distance="1350" swimtime="00:23:06.02" />
                    <SPLIT distance="1400" swimtime="00:23:58.18" />
                    <SPLIT distance="1450" swimtime="00:24:49.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="232" swimtime="00:03:25.17" resultid="9345" heatid="10714" lane="4" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                    <SPLIT distance="100" swimtime="00:01:38.09" />
                    <SPLIT distance="150" swimtime="00:02:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="205" swimtime="00:00:45.86" resultid="9346" heatid="10736" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1437" points="203" swimtime="00:01:38.73" resultid="9347" heatid="10840" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="9348" heatid="10874" lane="0" entrytime="00:07:15.00" />
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="9349" heatid="10895" lane="7" entrytime="00:03:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-03-21" firstname="Dariusz" gender="M" lastname="Wolny" nation="POL" athleteid="9339">
              <RESULTS>
                <RESULT eventid="1098" points="355" swimtime="00:10:37.95" resultid="9340" heatid="10673" lane="9" entrytime="00:10:22.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:01:15.76" />
                    <SPLIT distance="150" swimtime="00:01:53.54" />
                    <SPLIT distance="200" swimtime="00:02:32.22" />
                    <SPLIT distance="250" swimtime="00:03:10.92" />
                    <SPLIT distance="300" swimtime="00:03:50.23" />
                    <SPLIT distance="350" swimtime="00:04:29.81" />
                    <SPLIT distance="400" swimtime="00:05:09.68" />
                    <SPLIT distance="450" swimtime="00:05:49.62" />
                    <SPLIT distance="500" swimtime="00:06:30.17" />
                    <SPLIT distance="550" swimtime="00:07:10.98" />
                    <SPLIT distance="600" swimtime="00:07:52.14" />
                    <SPLIT distance="650" swimtime="00:08:33.38" />
                    <SPLIT distance="700" swimtime="00:09:15.30" />
                    <SPLIT distance="750" swimtime="00:09:57.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="373" swimtime="00:02:38.26" resultid="9341" heatid="10728" lane="4" entrytime="00:02:33.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:12.59" />
                    <SPLIT distance="150" swimtime="00:02:00.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="9342" heatid="10748" lane="5" entrytime="00:00:33.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-25" firstname="Marlena" gender="F" lastname="Jakubów" nation="POL" athleteid="9357">
              <RESULTS>
                <RESULT eventid="1059" points="192" swimtime="00:13:59.86" resultid="9358" heatid="10666" lane="4" entrytime="00:14:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.62" />
                    <SPLIT distance="100" swimtime="00:02:24.66" />
                    <SPLIT distance="150" swimtime="00:02:30.05" />
                    <SPLIT distance="250" swimtime="00:04:17.21" />
                    <SPLIT distance="350" swimtime="00:06:04.18" />
                    <SPLIT distance="450" swimtime="00:07:49.44" />
                    <SPLIT distance="550" swimtime="00:09:37.68" />
                    <SPLIT distance="650" swimtime="00:11:26.23" />
                    <SPLIT distance="750" swimtime="00:13:11.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="217" swimtime="00:00:45.03" resultid="9359" heatid="10736" lane="2" entrytime="00:00:44.00" />
                <RESULT eventid="1287" points="235" swimtime="00:01:24.35" resultid="9360" heatid="10768" lane="9" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="163" swimtime="00:01:46.30" resultid="9361" heatid="10840" lane="2" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="199" swimtime="00:03:13.51" resultid="9362" heatid="10852" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                    <SPLIT distance="100" swimtime="00:01:34.94" />
                    <SPLIT distance="150" swimtime="00:02:27.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="151" swimtime="00:03:52.78" resultid="9363" heatid="10895" lane="8" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.17" />
                    <SPLIT distance="100" swimtime="00:01:52.46" />
                    <SPLIT distance="150" swimtime="00:02:53.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="198" swimtime="00:06:45.67" resultid="9364" heatid="10931" lane="6" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                    <SPLIT distance="100" swimtime="00:01:33.44" />
                    <SPLIT distance="150" swimtime="00:02:26.30" />
                    <SPLIT distance="200" swimtime="00:03:19.92" />
                    <SPLIT distance="250" swimtime="00:04:12.97" />
                    <SPLIT distance="300" swimtime="00:05:05.36" />
                    <SPLIT distance="350" swimtime="00:05:58.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="260" swimtime="00:00:37.14" resultid="9804" heatid="10684" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1175" points="192" swimtime="00:03:38.39" resultid="9805" heatid="10714" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.71" />
                    <SPLIT distance="100" swimtime="00:01:49.13" />
                    <SPLIT distance="150" swimtime="00:02:52.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SPRZE" nation="POL" region="PDK" clubid="3424" name="GB Sport Rzeszów">
          <CONTACT email="marioss77rz@gmail.com" name="Mariusz Wójcicki" phone="660545998" />
          <ATHLETES>
            <ATHLETE birthdate="1973-09-05" firstname="Bartłomiej" gender="M" lastname="Czarnota" nation="POL" athleteid="3425">
              <RESULTS>
                <RESULT eventid="1098" points="333" swimtime="00:10:51.67" resultid="8005" heatid="10671" lane="6" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:12.06" />
                    <SPLIT distance="150" swimtime="00:01:52.25" />
                    <SPLIT distance="200" swimtime="00:02:33.12" />
                    <SPLIT distance="250" swimtime="00:03:14.14" />
                    <SPLIT distance="300" swimtime="00:03:55.43" />
                    <SPLIT distance="350" swimtime="00:04:36.91" />
                    <SPLIT distance="400" swimtime="00:05:18.46" />
                    <SPLIT distance="450" swimtime="00:05:59.22" />
                    <SPLIT distance="500" swimtime="00:06:40.58" />
                    <SPLIT distance="550" swimtime="00:07:22.59" />
                    <SPLIT distance="600" swimtime="00:08:05.08" />
                    <SPLIT distance="650" swimtime="00:08:46.75" />
                    <SPLIT distance="700" swimtime="00:09:29.37" />
                    <SPLIT distance="750" swimtime="00:10:12.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="494" swimtime="00:00:26.45" resultid="8006" heatid="10704" lane="3" entrytime="00:00:28.40" />
                <RESULT eventid="1272" points="421" swimtime="00:02:49.34" resultid="8007" heatid="10761" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:21.36" />
                    <SPLIT distance="150" swimtime="00:02:05.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="436" swimtime="00:01:15.29" resultid="8008" heatid="10815" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="8009" heatid="10863" lane="7" entrytime="00:02:20.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="8010" heatid="10920" lane="6" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-07-15" firstname="Grzegorz" gender="M" lastname="Wójcicki" nation="POL" athleteid="3432">
              <RESULTS>
                <RESULT eventid="1160" points="356" swimtime="00:00:29.49" resultid="8011" heatid="10704" lane="1" entrytime="00:00:28.60" />
                <RESULT eventid="1242" points="266" swimtime="00:00:37.35" resultid="8012" heatid="10746" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1302" points="314" swimtime="00:01:09.01" resultid="8013" heatid="10780" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="333" swimtime="00:00:32.33" resultid="8014" heatid="10832" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1638" points="291" swimtime="00:00:39.84" resultid="8015" heatid="10919" lane="2" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-11-19" firstname="Magdalena" gender="F" lastname="Jastrzębska" nation="POL" athleteid="3450">
              <RESULTS>
                <RESULT eventid="1226" points="97" swimtime="00:00:58.88" resultid="8026" heatid="10734" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="1376" points="189" swimtime="00:01:52.05" resultid="8027" heatid="10804" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="199" swimtime="00:00:50.43" resultid="8028" heatid="10906" lane="4" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-31" firstname="Sylwester" gender="M" lastname="Szewc" nation="POL" athleteid="3438">
              <RESULTS>
                <RESULT eventid="1160" points="394" swimtime="00:00:28.50" resultid="8016" heatid="10705" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1242" points="327" swimtime="00:00:34.86" resultid="8017" heatid="10747" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="359" swimtime="00:01:05.97" resultid="8018" heatid="10780" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="375" swimtime="00:00:31.09" resultid="8019" heatid="10831" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1638" points="292" swimtime="00:00:39.81" resultid="8020" heatid="10920" lane="7" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-01" firstname="Mariusz" gender="M" lastname="Wójcicki" nation="POL" athleteid="3444">
              <RESULTS>
                <RESULT eventid="1190" points="285" swimtime="00:02:53.15" resultid="8021" heatid="10724" lane="2" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:02:11.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="268" swimtime="00:02:52.89" resultid="8022" heatid="10795" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:18.62" />
                    <SPLIT distance="150" swimtime="00:02:05.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="288" swimtime="00:01:18.43" resultid="8023" heatid="10847" lane="5" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="242" swimtime="00:06:30.84" resultid="8024" heatid="10879" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="250" swimtime="00:03:57.86" />
                    <SPLIT distance="300" swimtime="00:04:57.36" />
                    <SPLIT distance="350" swimtime="00:05:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="326" swimtime="00:01:12.32" resultid="8025" heatid="10889" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="384" swimtime="00:02:08.49" resultid="8029" heatid="10802" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="150" swimtime="00:01:39.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3438" number="1" />
                    <RELAYPOSITION athleteid="3425" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3444" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3432" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" points="440" swimtime="00:01:51.52" resultid="8030" heatid="10872" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                    <SPLIT distance="100" swimtime="00:00:56.35" />
                    <SPLIT distance="150" swimtime="00:01:24.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3444" number="1" />
                    <RELAYPOSITION athleteid="3438" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3432" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3425" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAGDY" nation="POL" region="POM" clubid="9053" name="Gdynia Masters">
          <CONTACT email="k.mysiak@wpit.am.gdynia.pl" name="Mysiak" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Grażyna" gender="F" lastname="Heisler" nation="POL" athleteid="9067">
              <RESULTS>
                <RESULT eventid="1144" points="138" swimtime="00:00:45.91" resultid="9068" heatid="10681" lane="4" entrytime="00:00:49.00" />
                <RESULT eventid="1226" points="108" swimtime="00:00:56.66" resultid="9069" heatid="10735" lane="1" entrytime="00:00:56.00" />
                <RESULT eventid="1376" points="109" swimtime="00:02:14.33" resultid="9070" heatid="10803" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="117" swimtime="00:01:00.11" resultid="9071" heatid="10906" lane="2" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="9059">
              <RESULTS>
                <RESULT eventid="1160" points="154" swimtime="00:00:38.98" resultid="9060" heatid="10692" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1190" points="91" swimtime="00:04:13.34" resultid="9061" heatid="10720" lane="1" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.48" />
                    <SPLIT distance="100" swimtime="00:02:09.84" />
                    <SPLIT distance="150" swimtime="00:03:18.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="105" swimtime="00:00:50.86" resultid="9062" heatid="10743" lane="0" entrytime="00:00:50.00" />
                <RESULT eventid="1272" points="115" swimtime="00:04:20.91" resultid="9063" heatid="10758" lane="1" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.86" />
                    <SPLIT distance="100" swimtime="00:02:03.99" />
                    <SPLIT distance="150" swimtime="00:03:14.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="124" swimtime="00:01:54.32" resultid="9064" heatid="10811" lane="1" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="79" swimtime="00:02:00.61" resultid="9065" heatid="10844" lane="4" entrytime="00:01:58.00" />
                <RESULT eventid="1638" points="177" swimtime="00:00:46.97" resultid="9066" heatid="10915" lane="1" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="9072">
              <RESULTS>
                <RESULT eventid="1272" points="231" swimtime="00:03:26.91" resultid="9073" heatid="10759" lane="5" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.72" />
                    <SPLIT distance="100" swimtime="00:01:39.00" />
                    <SPLIT distance="150" swimtime="00:02:32.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="237" swimtime="00:01:32.28" resultid="9074" heatid="10813" lane="2" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="264" swimtime="00:00:41.14" resultid="9075" heatid="10917" lane="7" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Jan Maciej" gender="M" lastname="Boboli" nation="POL" athleteid="9054">
              <RESULTS>
                <RESULT eventid="1160" points="183" swimtime="00:00:36.83" resultid="9055" heatid="10693" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1242" points="67" swimtime="00:00:59.08" resultid="9056" heatid="10741" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1302" points="118" swimtime="00:01:35.63" resultid="9057" heatid="10774" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="154" swimtime="00:00:41.78" resultid="9058" heatid="10828" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="Ciundziewicki" nation="POL" athleteid="9076">
              <RESULTS>
                <RESULT eventid="1242" points="90" swimtime="00:00:53.46" resultid="9077" heatid="10741" lane="6" entrytime="00:00:57.00" />
                <RESULT eventid="1392" points="89" swimtime="00:02:07.76" resultid="9078" heatid="10810" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="69" swimtime="00:02:05.94" resultid="9079" heatid="10844" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="104" swimtime="00:00:56.03" resultid="9080" heatid="10914" lane="8" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="150" swimtime="00:02:55.54" resultid="9081" heatid="10800" lane="8" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.16" />
                    <SPLIT distance="150" swimtime="00:01:12.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9076" number="1" />
                    <RELAYPOSITION athleteid="9072" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9054" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9059" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" points="116" swimtime="00:02:53.53" resultid="9082" heatid="10870" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:01:39.58" />
                    <SPLIT distance="150" swimtime="00:02:15.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9059" number="1" />
                    <RELAYPOSITION athleteid="9076" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9072" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9054" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03714" nation="POL" region="14" clubid="9781" name="IKS Konstancin">
          <CONTACT email="plywalnia@ckr.pl" name="golon" />
          <ATHLETES>
            <ATHLETE birthdate="1971-02-23" firstname="Maciej" gender="M" lastname="Piłatowicz" nation="POL" athleteid="9782">
              <RESULTS>
                <RESULT eventid="1128" points="221" swimtime="00:23:59.93" resultid="9783" heatid="10676" lane="4" entrytime="00:24:30.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:24.54" />
                    <SPLIT distance="150" swimtime="00:02:11.10" />
                    <SPLIT distance="200" swimtime="00:02:57.66" />
                    <SPLIT distance="250" swimtime="00:03:45.83" />
                    <SPLIT distance="300" swimtime="00:04:33.91" />
                    <SPLIT distance="350" swimtime="00:05:21.49" />
                    <SPLIT distance="400" swimtime="00:06:10.01" />
                    <SPLIT distance="450" swimtime="00:06:57.85" />
                    <SPLIT distance="500" swimtime="00:07:45.96" />
                    <SPLIT distance="550" swimtime="00:08:34.72" />
                    <SPLIT distance="600" swimtime="00:09:22.95" />
                    <SPLIT distance="650" swimtime="00:10:12.02" />
                    <SPLIT distance="700" swimtime="00:11:01.31" />
                    <SPLIT distance="750" swimtime="00:11:49.96" />
                    <SPLIT distance="800" swimtime="00:12:38.36" />
                    <SPLIT distance="850" swimtime="00:13:26.95" />
                    <SPLIT distance="900" swimtime="00:14:15.79" />
                    <SPLIT distance="950" swimtime="00:15:04.71" />
                    <SPLIT distance="1000" swimtime="00:15:53.81" />
                    <SPLIT distance="1050" swimtime="00:16:42.64" />
                    <SPLIT distance="1100" swimtime="00:17:31.54" />
                    <SPLIT distance="1150" swimtime="00:18:19.32" />
                    <SPLIT distance="1200" swimtime="00:19:08.03" />
                    <SPLIT distance="1250" swimtime="00:19:57.10" />
                    <SPLIT distance="1300" swimtime="00:20:46.80" />
                    <SPLIT distance="1350" swimtime="00:21:35.64" />
                    <SPLIT distance="1400" swimtime="00:22:24.82" />
                    <SPLIT distance="1450" swimtime="00:23:13.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="9784" heatid="10831" lane="9" entrytime="00:00:33.11" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="9785" heatid="10888" lane="8" entrytime="00:01:18.11" />
                <RESULT eventid="1695" points="258" swimtime="00:05:45.60" resultid="9786" heatid="10940" lane="8" entrytime="00:05:55.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:02:01.24" />
                    <SPLIT distance="200" swimtime="00:02:45.75" />
                    <SPLIT distance="250" swimtime="00:03:30.88" />
                    <SPLIT distance="300" swimtime="00:04:16.01" />
                    <SPLIT distance="350" swimtime="00:05:01.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" region="14" clubid="3319" name="K.S.niezrzeszeni.pl">
          <CONTACT name="K.S.niezrzeszeni.pl" />
          <ATHLETES>
            <ATHLETE birthdate="1973-08-26" firstname="Małgorzata" gender="F" lastname="Piechura" nation="POL" athleteid="3336">
              <RESULTS>
                <RESULT eventid="1175" points="132" swimtime="00:04:07.61" resultid="6765" heatid="10713" lane="6" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.96" />
                    <SPLIT distance="100" swimtime="00:02:08.44" />
                    <SPLIT distance="150" swimtime="00:03:11.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="181" swimtime="00:04:05.76" resultid="6766" heatid="10754" lane="1" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.33" />
                    <SPLIT distance="100" swimtime="00:01:58.20" />
                    <SPLIT distance="150" swimtime="00:03:01.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="141" swimtime="00:03:37.01" resultid="6767" heatid="10852" lane="0" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.72" />
                    <SPLIT distance="100" swimtime="00:01:40.44" />
                    <SPLIT distance="150" swimtime="00:02:39.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="132" swimtime="00:07:44.31" resultid="6768" heatid="10931" lane="4" entrytime="00:07:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.07" />
                    <SPLIT distance="100" swimtime="00:01:45.37" />
                    <SPLIT distance="150" swimtime="00:02:44.44" />
                    <SPLIT distance="200" swimtime="00:03:43.58" />
                    <SPLIT distance="250" swimtime="00:04:44.03" />
                    <SPLIT distance="300" swimtime="00:05:46.68" />
                    <SPLIT distance="350" swimtime="00:06:49.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="3328">
              <RESULTS>
                <RESULT eventid="1128" points="193" swimtime="00:25:06.84" resultid="6758" heatid="10676" lane="3" entrytime="00:24:58.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.63" />
                    <SPLIT distance="100" swimtime="00:01:29.14" />
                    <SPLIT distance="150" swimtime="00:02:17.06" />
                    <SPLIT distance="200" swimtime="00:03:07.33" />
                    <SPLIT distance="250" swimtime="00:03:56.61" />
                    <SPLIT distance="300" swimtime="00:04:46.50" />
                    <SPLIT distance="350" swimtime="00:05:36.75" />
                    <SPLIT distance="400" swimtime="00:06:27.25" />
                    <SPLIT distance="450" swimtime="00:07:17.41" />
                    <SPLIT distance="500" swimtime="00:08:07.65" />
                    <SPLIT distance="550" swimtime="00:08:58.30" />
                    <SPLIT distance="600" swimtime="00:09:49.77" />
                    <SPLIT distance="650" swimtime="00:10:40.51" />
                    <SPLIT distance="700" swimtime="00:11:31.94" />
                    <SPLIT distance="750" swimtime="00:12:23.31" />
                    <SPLIT distance="800" swimtime="00:13:14.79" />
                    <SPLIT distance="850" swimtime="00:14:06.34" />
                    <SPLIT distance="900" swimtime="00:14:58.67" />
                    <SPLIT distance="950" swimtime="00:15:50.14" />
                    <SPLIT distance="1000" swimtime="00:16:42.63" />
                    <SPLIT distance="1050" swimtime="00:17:35.16" />
                    <SPLIT distance="1100" swimtime="00:18:26.77" />
                    <SPLIT distance="1150" swimtime="00:19:18.22" />
                    <SPLIT distance="1200" swimtime="00:20:10.54" />
                    <SPLIT distance="1250" swimtime="00:21:01.05" />
                    <SPLIT distance="1300" swimtime="00:21:51.61" />
                    <SPLIT distance="1350" swimtime="00:22:42.10" />
                    <SPLIT distance="1400" swimtime="00:23:33.27" />
                    <SPLIT distance="1450" swimtime="00:24:22.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="205" swimtime="00:00:35.45" resultid="6759" heatid="10690" lane="6" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="6760" heatid="10721" lane="6" entrytime="00:03:28.20" />
                <RESULT eventid="1242" points="195" swimtime="00:00:41.44" resultid="6761" heatid="10744" lane="5" entrytime="00:00:41.17" />
                <RESULT eventid="1302" points="212" swimtime="00:01:18.59" resultid="6762" heatid="10775" lane="3" entrytime="00:01:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="192" swimtime="00:01:29.87" resultid="6763" heatid="10846" lane="0" entrytime="00:01:31.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="193" swimtime="00:03:13.49" resultid="6764" heatid="10901" lane="7" entrytime="00:03:15.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                    <SPLIT distance="100" swimtime="00:01:34.42" />
                    <SPLIT distance="150" swimtime="00:02:25.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KATAK" nation="LTU" clubid="4651" name="Kauno Takas">
          <CONTACT city="Kaunas" email="kaunotakas@gmail.com" internet="klubastakas.lt" name="Linas Kersevicius" phone="+37068780249" street="Lentvario g. 19" zip="44439" />
          <ATHLETES>
            <ATHLETE birthdate="1969-08-22" firstname="Arvydas" gender="M" lastname="Burinskas" nation="LTU" athleteid="4662">
              <RESULTS>
                <RESULT eventid="1332" points="252" swimtime="00:02:56.49" resultid="8206" heatid="10794" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:22.83" />
                    <SPLIT distance="150" swimtime="00:02:09.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="389" swimtime="00:00:30.71" resultid="8207" heatid="10834" lane="7" entrytime="00:00:30.20" />
                <RESULT eventid="1578" points="286" swimtime="00:01:15.57" resultid="8208" heatid="10888" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-08" firstname="Pavelas" gender="M" lastname="Bezzubovas" nation="LTU" athleteid="4666">
              <RESULTS>
                <RESULT eventid="1160" points="169" swimtime="00:00:37.81" resultid="8209" heatid="10693" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1422" points="68" swimtime="00:00:54.80" resultid="8210" heatid="10827" lane="3" entrytime="00:00:44.00" />
                <RESULT eventid="1638" points="136" swimtime="00:00:51.29" resultid="8211" heatid="10914" lane="7" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-06-18" firstname="Linas" gender="M" lastname="Kersevicius" nation="LTU" athleteid="4652">
              <RESULTS>
                <RESULT eventid="1160" points="397" swimtime="00:00:28.44" resultid="8198" heatid="10702" lane="0" entrytime="00:00:29.50" />
                <RESULT eventid="1242" points="406" swimtime="00:00:32.44" resultid="8199" heatid="10749" lane="1" entrytime="00:00:32.50" />
                <RESULT eventid="1452" points="397" swimtime="00:01:10.52" resultid="8200" heatid="10849" lane="0" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="388" swimtime="00:02:33.40" resultid="8201" heatid="10903" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                    <SPLIT distance="100" swimtime="00:01:14.25" />
                    <SPLIT distance="150" swimtime="00:01:54.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-06" firstname="Vedestas" gender="M" lastname="Sefleris" nation="LTU" athleteid="4657">
              <RESULTS>
                <RESULT eventid="1332" points="402" swimtime="00:02:30.97" resultid="8202" heatid="10796" lane="8" entrytime="00:02:30.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:01:09.06" />
                    <SPLIT distance="150" swimtime="00:01:47.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="504" swimtime="00:00:28.18" resultid="8203" heatid="10836" lane="3" entrytime="00:00:28.35" />
                <RESULT eventid="1578" points="496" swimtime="00:01:02.93" resultid="8204" heatid="10891" lane="7" entrytime="00:01:04.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="8205" heatid="10942" lane="9" entrytime="00:05:20.10" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KSMAK" nation="POL" region="MAZ" clubid="4446" name="Klub Sportowy Mako">
          <CONTACT email="ania.plywanie@gmail.com" name="Anna Dąbrowska" phone="601480280" />
          <ATHLETES>
            <ATHLETE birthdate="1980-06-07" firstname="Piotr" gender="M" lastname="Kieżun" nation="POL" athleteid="4464">
              <RESULTS>
                <RESULT eventid="1160" points="269" swimtime="00:00:32.38" resultid="6997" heatid="10697" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1302" points="250" swimtime="00:01:14.41" resultid="6998" heatid="10778" lane="3" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="257" swimtime="00:00:41.51" resultid="6999" heatid="10918" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-20" firstname="Anna" gender="F" lastname="Dąbrowska" nation="POL" athleteid="4474">
              <RESULTS>
                <RESULT eventid="1144" points="265" swimtime="00:00:36.91" resultid="7004" heatid="10684" lane="5" entrytime="00:00:35.60" />
                <RESULT eventid="1287" points="245" swimtime="00:01:23.14" resultid="7005" heatid="10767" lane="4" entrytime="00:01:22.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="221" swimtime="00:00:40.39" resultid="7006" heatid="10821" lane="3" entrytime="00:00:42.30" />
                <RESULT eventid="1562" points="178" swimtime="00:01:38.53" resultid="7007" heatid="10883" lane="7" entrytime="00:01:41.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-06-01" firstname="Robert" gender="M" lastname="Wilk" nation="POL" athleteid="4484">
              <RESULTS>
                <RESULT eventid="1422" points="586" swimtime="00:00:26.79" resultid="7011" heatid="10838" lane="8" entrytime="00:00:26.17" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-07" firstname="Sławomir" gender="M" lastname="Szcześniak" nation="POL" athleteid="4499">
              <RESULTS>
                <RESULT eventid="1160" points="332" swimtime="00:00:30.17" resultid="7021" heatid="10696" lane="4" entrytime="00:00:33.50" />
                <RESULT eventid="1302" points="216" swimtime="00:01:18.17" resultid="7022" heatid="10775" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 15 - Brak dotknięcia ściany obydwiema rozłaczonymi dłońmi przy nawrocie lub na zakończenie wyścigu" eventid="1392" status="DSQ" swimtime="00:01:30.97" resultid="7023" heatid="10814" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="7024" heatid="10829" lane="2" entrytime="00:00:36.00" />
                <RESULT comment="K 15 - Brak dotknięcia ściany obydwiema rozłaczonymi dłońmi przy nawrocie lub na zakończenie wyścigu" eventid="1638" status="DSQ" swimtime="00:00:40.17" resultid="7025" heatid="10920" lane="9" entrytime="00:00:38.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-06-25" firstname="Krzysztof" gender="M" lastname="Wilk" nation="POL" athleteid="4486">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="7012" heatid="10711" lane="0" entrytime="00:00:24.70" />
                <RESULT eventid="1302" points="588" swimtime="00:00:55.98" resultid="7013" heatid="10788" lane="8" entrytime="00:00:55.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="7014" heatid="10866" lane="1" entrytime="00:02:07.07" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-05-14" firstname="Dominik" gender="M" lastname="Markowski" nation="POL" athleteid="4472">
              <RESULTS>
                <RESULT eventid="1695" points="163" swimtime="00:06:42.16" resultid="7003" heatid="10937" lane="6" entrytime="00:06:45.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                    <SPLIT distance="100" swimtime="00:01:34.12" />
                    <SPLIT distance="150" swimtime="00:02:25.70" />
                    <SPLIT distance="200" swimtime="00:03:17.41" />
                    <SPLIT distance="250" swimtime="00:04:09.56" />
                    <SPLIT distance="300" swimtime="00:05:02.10" />
                    <SPLIT distance="350" swimtime="00:05:55.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-20" firstname="Jacek" gender="M" lastname="Suda" nation="POL" athleteid="4494">
              <RESULTS>
                <RESULT eventid="1160" points="260" swimtime="00:00:32.75" resultid="7018" heatid="10696" lane="7" entrytime="00:00:34.70" />
                <RESULT eventid="1302" points="278" swimtime="00:01:11.81" resultid="7019" heatid="10777" lane="9" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-30" firstname="Piotr" gender="M" lastname="Safrończyk" nation="POL" athleteid="4479">
              <RESULTS>
                <RESULT eventid="1160" points="590" swimtime="00:00:24.93" resultid="7008" heatid="10710" lane="4" entrytime="00:00:24.90" />
                <RESULT eventid="1638" points="657" swimtime="00:00:30.39" resultid="7009" heatid="10926" lane="2" entrytime="00:00:30.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-13" firstname="Jacek" gender="M" lastname="Kalwasiński" nation="POL" athleteid="4497">
              <RESULTS>
                <RESULT comment="O 4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1160" status="DSQ" swimtime="00:00:32.65" resultid="7020" heatid="10698" lane="7" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-23" firstname="Katarzyna" gender="F" lastname="Żołnowska" nation="POL" athleteid="4505">
              <RESULTS>
                <RESULT eventid="1175" points="581" swimtime="00:02:31.07" resultid="7026" heatid="10718" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                    <SPLIT distance="150" swimtime="00:01:55.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-09" firstname="Paweł" gender="M" lastname="Rurak" nation="POL" athleteid="4461" />
            <ATHLETE birthdate="1978-04-07" firstname="Tomasz" gender="M" lastname="Jurkowski" nation="POL" athleteid="4468">
              <RESULTS>
                <RESULT eventid="1160" points="310" swimtime="00:00:30.87" resultid="7000" heatid="10696" lane="2" entrytime="00:00:34.73" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="7001" heatid="10721" lane="2" entrytime="00:03:28.94" />
                <RESULT eventid="1638" points="289" swimtime="00:00:39.93" resultid="7002" heatid="10918" lane="6" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-29" firstname="Artur" gender="M" lastname="Pietrzak" nation="POL" athleteid="4482">
              <RESULTS>
                <RESULT eventid="1422" points="534" swimtime="00:00:27.64" resultid="7010" heatid="10835" lane="2" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  w  kat A  100-119  lat" eventid="1368" points="617" swimtime="00:01:49.71" resultid="7027" heatid="10802" lane="5" entrytime="00:01:52.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:00:57.93" />
                    <SPLIT distance="150" swimtime="00:01:25.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4461" number="1" />
                    <RELAYPOSITION athleteid="4479" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4482" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4486" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1368" points="195" swimtime="00:02:40.91" resultid="7029" heatid="10800" lane="3" entrytime="00:02:30.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:01:23.30" />
                    <SPLIT distance="150" swimtime="00:02:09.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4468" number="1" />
                    <RELAYPOSITION athleteid="4464" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4499" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4497" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn w  kat A  100-119  lat" eventid="1518" points="663" swimtime="00:01:37.27" resultid="7030" heatid="10872" lane="5" entrytime="00:01:38.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.74" />
                    <SPLIT distance="100" swimtime="00:00:48.69" />
                    <SPLIT distance="150" swimtime="00:01:12.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4484" number="1" />
                    <RELAYPOSITION athleteid="4479" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4461" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4486" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1518" points="286" swimtime="00:02:08.73" resultid="7031" heatid="10870" lane="2" entrytime="00:02:15.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:04.60" />
                    <SPLIT distance="150" swimtime="00:01:36.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4464" number="1" />
                    <RELAYPOSITION athleteid="4468" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4494" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4499" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:01:54.10" resultid="7028" heatid="10733" lane="2" entrytime="00:01:54.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.74" />
                    <SPLIT distance="100" swimtime="00:00:53.29" />
                    <SPLIT distance="150" swimtime="00:01:30.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4479" number="1" />
                    <RELAYPOSITION athleteid="4505" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4474" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4486" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:05.81" resultid="7032" heatid="10929" lane="1" entrytime="00:02:09.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4461" number="1" />
                    <RELAYPOSITION athleteid="4479" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4505" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4474" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WAPOZ" nation="POL" region="WIE" clubid="5973" name="Klub Sportowy Warta Poznań">
          <CONTACT city="Poznań" email="jacek.thiem@gmail.com" name="Jacek Thiem" phone="502499565" state="WIE" street="Osiedle Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1957-10-01" firstname="Rusłana" gender="F" lastname="Dembecka" nation="POL" license="100115600353" athleteid="9601">
              <RESULTS>
                <RESULT eventid="1059" points="69" swimtime="00:19:38.64" resultid="9602" heatid="10666" lane="0" entrytime="00:18:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.68" />
                    <SPLIT distance="100" swimtime="00:02:07.62" />
                    <SPLIT distance="150" swimtime="00:03:23.05" />
                    <SPLIT distance="200" swimtime="00:04:40.90" />
                    <SPLIT distance="250" swimtime="00:05:57.43" />
                    <SPLIT distance="300" swimtime="00:07:16.63" />
                    <SPLIT distance="350" swimtime="00:08:32.81" />
                    <SPLIT distance="400" swimtime="00:09:48.19" />
                    <SPLIT distance="450" swimtime="00:11:03.84" />
                    <SPLIT distance="500" swimtime="00:12:18.75" />
                    <SPLIT distance="550" swimtime="00:13:33.21" />
                    <SPLIT distance="600" swimtime="00:14:48.83" />
                    <SPLIT distance="650" swimtime="00:16:01.90" />
                    <SPLIT distance="700" swimtime="00:17:15.32" />
                    <SPLIT distance="750" swimtime="00:18:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="98" swimtime="00:00:51.45" resultid="9603" heatid="10682" lane="9" entrytime="00:00:49.00" />
                <RESULT eventid="1226" points="71" swimtime="00:01:05.15" resultid="9604" heatid="10734" lane="6" entrytime="00:01:04.00" />
                <RESULT eventid="1257" points="144" swimtime="00:04:25.22" resultid="9605" heatid="10753" lane="2" entrytime="00:04:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.62" />
                    <SPLIT distance="100" swimtime="00:02:08.65" />
                    <SPLIT distance="150" swimtime="00:03:18.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="133" swimtime="00:02:05.95" resultid="9606" heatid="10804" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="73" swimtime="00:04:30.25" resultid="9607" heatid="10851" lane="2" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.27" />
                    <SPLIT distance="100" swimtime="00:02:08.63" />
                    <SPLIT distance="150" swimtime="00:03:20.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="52" swimtime="00:05:30.54" resultid="9608" heatid="10894" lane="0" entrytime="00:04:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.14" />
                    <SPLIT distance="100" swimtime="00:02:44.38" />
                    <SPLIT distance="150" swimtime="00:04:12.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="75" swimtime="00:09:19.76" resultid="9609" heatid="10931" lane="9" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.14" />
                    <SPLIT distance="100" swimtime="00:02:06.88" />
                    <SPLIT distance="150" swimtime="00:03:18.81" />
                    <SPLIT distance="200" swimtime="00:04:31.43" />
                    <SPLIT distance="250" swimtime="00:05:45.47" />
                    <SPLIT distance="300" swimtime="00:06:57.95" />
                    <SPLIT distance="350" swimtime="00:08:10.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="Kaczmarek" nation="POL" license="100115700354" athleteid="9582">
              <RESULTS>
                <RESULT eventid="1098" points="517" swimtime="00:09:23.26" resultid="9583" heatid="10673" lane="5" entrytime="00:09:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:43.24" />
                    <SPLIT distance="200" swimtime="00:02:19.64" />
                    <SPLIT distance="250" swimtime="00:02:55.45" />
                    <SPLIT distance="300" swimtime="00:03:31.30" />
                    <SPLIT distance="350" swimtime="00:04:06.86" />
                    <SPLIT distance="400" swimtime="00:04:41.56" />
                    <SPLIT distance="450" swimtime="00:05:16.58" />
                    <SPLIT distance="500" swimtime="00:05:52.08" />
                    <SPLIT distance="550" swimtime="00:06:27.33" />
                    <SPLIT distance="600" swimtime="00:07:03.11" />
                    <SPLIT distance="650" swimtime="00:07:38.65" />
                    <SPLIT distance="700" swimtime="00:08:14.25" />
                    <SPLIT distance="750" swimtime="00:08:49.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="511" swimtime="00:02:22.51" resultid="9584" heatid="10730" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                    <SPLIT distance="100" swimtime="00:01:08.36" />
                    <SPLIT distance="150" swimtime="00:01:49.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="473" swimtime="00:02:42.91" resultid="9585" heatid="10764" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                    <SPLIT distance="100" swimtime="00:01:18.11" />
                    <SPLIT distance="150" swimtime="00:02:00.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="482" swimtime="00:02:22.22" resultid="9586" heatid="10796" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:08.43" />
                    <SPLIT distance="150" swimtime="00:01:44.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="504" swimtime="00:02:08.16" resultid="9587" heatid="10866" lane="6" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:05.02" />
                    <SPLIT distance="150" swimtime="00:01:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="483" swimtime="00:05:10.65" resultid="9588" heatid="10881" lane="6" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:07.81" />
                    <SPLIT distance="150" swimtime="00:01:52.40" />
                    <SPLIT distance="200" swimtime="00:02:34.68" />
                    <SPLIT distance="250" swimtime="00:03:18.51" />
                    <SPLIT distance="300" swimtime="00:04:02.70" />
                    <SPLIT distance="350" swimtime="00:04:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="475" swimtime="00:01:03.82" resultid="9589" heatid="10891" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="518" swimtime="00:04:34.02" resultid="9590" heatid="10945" lane="5" entrytime="00:04:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:06.41" />
                    <SPLIT distance="150" swimtime="00:01:41.47" />
                    <SPLIT distance="200" swimtime="00:02:17.10" />
                    <SPLIT distance="250" swimtime="00:02:51.71" />
                    <SPLIT distance="300" swimtime="00:03:26.52" />
                    <SPLIT distance="350" swimtime="00:04:00.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-02" firstname="Tomasz" gender="M" lastname="Tomaszewski" nation="POL" license="500115700466" athleteid="9628">
              <RESULTS>
                <RESULT eventid="1242" points="465" swimtime="00:00:31.01" resultid="9629" heatid="10750" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1452" points="462" swimtime="00:01:07.03" resultid="9630" heatid="10849" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="9631" heatid="10862" lane="8" entrytime="00:02:28.00" />
                <RESULT eventid="1608" points="402" swimtime="00:02:31.58" resultid="9632" heatid="10903" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:14.11" />
                    <SPLIT distance="150" swimtime="00:01:54.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-03" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" license="100115700350" athleteid="9618">
              <RESULTS>
                <RESULT eventid="1160" points="405" swimtime="00:00:28.25" resultid="9619" heatid="10703" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1302" points="442" swimtime="00:01:01.56" resultid="9620" heatid="10783" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="366" swimtime="00:00:31.33" resultid="9621" heatid="10832" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1695" points="397" swimtime="00:04:59.30" resultid="9622" heatid="10943" lane="9" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                    <SPLIT distance="150" swimtime="00:01:50.43" />
                    <SPLIT distance="200" swimtime="00:02:29.03" />
                    <SPLIT distance="250" swimtime="00:03:07.62" />
                    <SPLIT distance="300" swimtime="00:03:46.26" />
                    <SPLIT distance="350" swimtime="00:04:23.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-31" firstname="Bartłomiej" gender="M" lastname="Zadorożny" nation="POL" license="500115700461" athleteid="9610">
              <RESULTS>
                <RESULT eventid="1160" points="429" swimtime="00:00:27.72" resultid="9611" heatid="10705" lane="3" entrytime="00:00:27.74" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="9612" heatid="10725" lane="4" entrytime="00:02:47.06" />
                <RESULT eventid="1272" points="392" swimtime="00:02:53.49" resultid="9613" heatid="10762" lane="4" entrytime="00:02:53.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:19.87" />
                    <SPLIT distance="150" swimtime="00:02:04.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="381" swimtime="00:01:04.69" resultid="9614" heatid="10784" lane="9" entrytime="00:01:02.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="445" swimtime="00:01:14.79" resultid="9615" heatid="10817" lane="4" entrytime="00:01:16.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="357" swimtime="00:00:31.61" resultid="9616" heatid="10833" lane="1" entrytime="00:00:30.98" />
                <RESULT eventid="1638" points="491" swimtime="00:00:33.47" resultid="9617" heatid="10924" lane="0" entrytime="00:00:34.16" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-07-13" firstname="Paulina" gender="F" lastname="Mendowska" nation="POL" athleteid="9633">
              <RESULTS>
                <RESULT eventid="1376" points="417" swimtime="00:01:26.08" resultid="9634" heatid="10808" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="428" swimtime="00:00:32.40" resultid="9635" heatid="10824" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1562" points="472" swimtime="00:01:11.21" resultid="9636" heatid="10884" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="425" swimtime="00:02:45.00" resultid="9637" heatid="10897" lane="4" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:20.65" />
                    <SPLIT distance="150" swimtime="00:02:03.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-10-01" firstname="Grażyna" gender="F" lastname="Drela" nation="POL" license="500115700493" athleteid="9577">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat H  60-64 lat" eventid="1175" points="280" swimtime="00:03:12.73" resultid="9578" heatid="10714" lane="6" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:30.57" />
                    <SPLIT distance="150" swimtime="00:02:24.41" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat H  60-64 lata" eventid="1257" points="296" swimtime="00:03:28.61" resultid="9579" heatid="10755" lane="8" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.86" />
                    <SPLIT distance="100" swimtime="00:01:41.26" />
                    <SPLIT distance="150" swimtime="00:02:37.20" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat H  60-64  lat" eventid="1376" points="318" swimtime="00:01:34.26" resultid="9580" heatid="10806" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1623" points="318" swimtime="00:00:43.18" resultid="9581" heatid="10909" lane="9" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="Waraczewski" nation="POL" license="100115700344" athleteid="9623">
              <RESULTS>
                <RESULT eventid="1190" points="238" swimtime="00:03:03.73" resultid="9624" heatid="10723" lane="1" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:01:31.44" />
                    <SPLIT distance="150" swimtime="00:02:23.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="289" swimtime="00:03:12.01" resultid="9625" heatid="10761" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:01:31.60" />
                    <SPLIT distance="150" swimtime="00:02:23.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="280" swimtime="00:01:27.27" resultid="9626" heatid="10814" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="305" swimtime="00:00:39.21" resultid="9627" heatid="10918" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-08" firstname="Katarzyna" gender="F" lastname="Mendowska" nation="POL" athleteid="9638">
              <RESULTS>
                <RESULT comment="M 1 - Głowa pływaka nie złamała lustra wody przed lub na linii 15 m" eventid="1562" status="DSQ" swimtime="00:01:13.30" resultid="9639" heatid="10884" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="451" swimtime="00:02:41.72" resultid="9640" heatid="10897" lane="5" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                    <SPLIT distance="100" swimtime="00:01:19.65" />
                    <SPLIT distance="150" swimtime="00:02:01.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-22" firstname="Małgorzata" gender="F" lastname="Putowska" nation="POL" license="500115600462" athleteid="9591">
              <RESULTS>
                <RESULT eventid="1059" points="128" swimtime="00:16:00.29" resultid="9592" heatid="10666" lane="2" entrytime="00:16:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                    <SPLIT distance="100" swimtime="00:01:45.14" />
                    <SPLIT distance="150" swimtime="00:02:44.89" />
                    <SPLIT distance="200" swimtime="00:03:46.58" />
                    <SPLIT distance="250" swimtime="00:04:49.26" />
                    <SPLIT distance="300" swimtime="00:05:51.13" />
                    <SPLIT distance="350" swimtime="00:06:54.03" />
                    <SPLIT distance="400" swimtime="00:07:56.07" />
                    <SPLIT distance="450" swimtime="00:08:58.15" />
                    <SPLIT distance="500" swimtime="00:09:59.16" />
                    <SPLIT distance="550" swimtime="00:11:00.89" />
                    <SPLIT distance="600" swimtime="00:12:01.70" />
                    <SPLIT distance="650" swimtime="00:13:02.03" />
                    <SPLIT distance="700" swimtime="00:14:02.65" />
                    <SPLIT distance="750" swimtime="00:15:02.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="199" swimtime="00:00:40.60" resultid="9593" heatid="10682" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1175" points="143" swimtime="00:04:00.62" resultid="9594" heatid="10714" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.89" />
                    <SPLIT distance="100" swimtime="00:01:58.45" />
                    <SPLIT distance="150" swimtime="00:03:06.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="173" swimtime="00:04:09.20" resultid="9595" heatid="10754" lane="8" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.48" />
                    <SPLIT distance="100" swimtime="00:02:00.75" />
                    <SPLIT distance="150" swimtime="00:03:07.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1317" points="74" swimtime="00:04:49.29" resultid="9596" heatid="10790" lane="9" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.16" />
                    <SPLIT distance="100" swimtime="00:02:15.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="124" swimtime="00:01:56.38" resultid="9597" heatid="10840" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="144" swimtime="00:08:27.11" resultid="9598" heatid="10873" lane="4" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.78" />
                    <SPLIT distance="100" swimtime="00:02:10.89" />
                    <SPLIT distance="150" swimtime="00:03:13.62" />
                    <SPLIT distance="200" swimtime="00:04:15.93" />
                    <SPLIT distance="250" swimtime="00:05:23.67" />
                    <SPLIT distance="300" swimtime="00:06:29.94" />
                    <SPLIT distance="350" swimtime="00:07:26.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="73" swimtime="00:02:12.39" resultid="9599" heatid="10883" lane="0" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="124" swimtime="00:04:08.51" resultid="9600" heatid="10894" lane="5" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.94" />
                    <SPLIT distance="100" swimtime="00:02:01.07" />
                    <SPLIT distance="150" swimtime="00:03:05.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1368" points="462" swimtime="00:02:00.84" resultid="9642" heatid="10801" lane="4" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:01:04.37" />
                    <SPLIT distance="150" swimtime="00:01:32.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9628" number="1" />
                    <RELAYPOSITION athleteid="9610" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9582" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9618" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1518" points="391" swimtime="00:01:55.94" resultid="9643" heatid="10871" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                    <SPLIT distance="100" swimtime="00:00:54.71" />
                    <SPLIT distance="150" swimtime="00:01:27.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9628" number="1" />
                    <RELAYPOSITION athleteid="9610" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9623" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9618" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:15.86" resultid="9641" heatid="10732" lane="9" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                    <SPLIT distance="100" swimtime="00:01:02.55" />
                    <SPLIT distance="150" swimtime="00:02:00.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9628" number="1" />
                    <RELAYPOSITION athleteid="9577" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9591" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9623" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:39.06" resultid="9644" heatid="10928" lane="7" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:02:05.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9628" number="1" />
                    <RELAYPOSITION athleteid="9577" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9591" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9623" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KOKRA" nation="POL" region="MAL" clubid="4150" name="Korona Kraków Masters">
          <CONTACT city="Kraków" name="Mariola Kuliś" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1982-02-08" firstname="Tomasz" gender="M" lastname="Czerniecki" nation="POL" athleteid="4216">
              <RESULTS>
                <RESULT eventid="1160" points="520" swimtime="00:00:25.99" resultid="6658" heatid="10709" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1302" points="486" swimtime="00:00:59.66" resultid="6659" heatid="10786" lane="4" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="6660" heatid="10835" lane="3" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="4203">
              <RESULTS>
                <RESULT eventid="1175" points="300" swimtime="00:03:08.33" resultid="6648" heatid="10715" lane="5" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                    <SPLIT distance="100" swimtime="00:01:28.38" />
                    <SPLIT distance="150" swimtime="00:02:24.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="283" swimtime="00:06:45.54" resultid="6649" heatid="10874" lane="6" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:28.01" />
                    <SPLIT distance="150" swimtime="00:02:24.94" />
                    <SPLIT distance="200" swimtime="00:03:19.52" />
                    <SPLIT distance="250" swimtime="00:04:17.60" />
                    <SPLIT distance="300" swimtime="00:05:15.70" />
                    <SPLIT distance="350" swimtime="00:06:02.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="265" swimtime="00:01:26.32" resultid="6650" heatid="10884" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="4151">
              <RESULTS>
                <RESULT eventid="1144" points="486" swimtime="00:00:30.17" resultid="6604" heatid="10687" lane="4" entrytime="00:00:29.85" />
                <RESULT eventid="1226" points="401" swimtime="00:00:36.69" resultid="6605" heatid="10738" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1287" points="423" swimtime="00:01:09.31" resultid="6606" heatid="10770" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="403" swimtime="00:00:33.05" resultid="6607" heatid="10822" lane="2" entrytime="00:00:38.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat F  50-54  lata" eventid="1437" points="368" swimtime="00:01:21.07" resultid="6608" heatid="10842" lane="0" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="472" swimtime="00:00:37.84" resultid="6609" heatid="10911" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-29" firstname="Jolanta" gender="F" lastname="Uczarczyk" nation="POL" athleteid="4190">
              <RESULTS>
                <RESULT eventid="1144" points="245" swimtime="00:00:37.90" resultid="6637" heatid="10683" lane="3" entrytime="00:00:38.48" />
                <RESULT eventid="1175" points="161" swimtime="00:03:51.44" resultid="6638" heatid="10713" lane="3" entrytime="00:03:52.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="100" swimtime="00:01:49.02" />
                    <SPLIT distance="150" swimtime="00:02:57.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="161" swimtime="00:00:49.67" resultid="6639" heatid="10736" lane="3" entrytime="00:00:43.00" />
                <RESULT eventid="1287" points="196" swimtime="00:01:29.60" resultid="6640" heatid="10767" lane="7" entrytime="00:01:27.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="167" swimtime="00:00:44.29" resultid="6641" heatid="10821" lane="7" entrytime="00:00:46.36" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-30" firstname="Piotr" gender="M" lastname="Łysiak" nation="POL" athleteid="4158">
              <RESULTS>
                <RESULT eventid="1272" points="363" swimtime="00:02:57.97" resultid="6610" heatid="10762" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:22.42" />
                    <SPLIT distance="150" swimtime="00:02:07.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="337" swimtime="00:01:22.07" resultid="6611" heatid="10816" lane="8" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="352" swimtime="00:00:37.39" resultid="6612" heatid="10922" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-12-18" firstname="Szymon" gender="M" lastname="Pyrć" nation="POL" athleteid="4187">
              <RESULTS>
                <RESULT eventid="1128" points="372" swimtime="00:20:10.77" resultid="6635" heatid="10679" lane="9" entrytime="00:20:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:01:56.57" />
                    <SPLIT distance="200" swimtime="00:02:37.40" />
                    <SPLIT distance="250" swimtime="00:03:18.22" />
                    <SPLIT distance="300" swimtime="00:03:59.26" />
                    <SPLIT distance="350" swimtime="00:04:40.10" />
                    <SPLIT distance="400" swimtime="00:05:20.88" />
                    <SPLIT distance="450" swimtime="00:06:01.50" />
                    <SPLIT distance="500" swimtime="00:06:42.19" />
                    <SPLIT distance="550" swimtime="00:07:23.13" />
                    <SPLIT distance="600" swimtime="00:08:03.65" />
                    <SPLIT distance="650" swimtime="00:08:44.67" />
                    <SPLIT distance="700" swimtime="00:09:25.08" />
                    <SPLIT distance="750" swimtime="00:10:05.53" />
                    <SPLIT distance="800" swimtime="00:10:45.90" />
                    <SPLIT distance="850" swimtime="00:11:26.28" />
                    <SPLIT distance="900" swimtime="00:12:06.51" />
                    <SPLIT distance="950" swimtime="00:12:47.37" />
                    <SPLIT distance="1000" swimtime="00:13:27.93" />
                    <SPLIT distance="1050" swimtime="00:14:08.68" />
                    <SPLIT distance="1100" swimtime="00:14:49.15" />
                    <SPLIT distance="1150" swimtime="00:15:29.69" />
                    <SPLIT distance="1200" swimtime="00:16:10.31" />
                    <SPLIT distance="1250" swimtime="00:16:50.84" />
                    <SPLIT distance="1300" swimtime="00:17:31.44" />
                    <SPLIT distance="1350" swimtime="00:18:11.84" />
                    <SPLIT distance="1400" swimtime="00:18:52.38" />
                    <SPLIT distance="1450" swimtime="00:19:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="367" swimtime="00:02:35.71" resultid="6636" heatid="10795" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:12.20" />
                    <SPLIT distance="150" swimtime="00:01:52.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="4220">
              <RESULTS>
                <RESULT eventid="1059" points="255" swimtime="00:12:44.48" resultid="6661" heatid="10667" lane="2" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                    <SPLIT distance="100" swimtime="00:01:25.71" />
                    <SPLIT distance="150" swimtime="00:02:13.08" />
                    <SPLIT distance="200" swimtime="00:03:00.12" />
                    <SPLIT distance="250" swimtime="00:03:48.28" />
                    <SPLIT distance="300" swimtime="00:04:37.86" />
                    <SPLIT distance="350" swimtime="00:05:27.23" />
                    <SPLIT distance="400" swimtime="00:06:16.83" />
                    <SPLIT distance="450" swimtime="00:07:06.49" />
                    <SPLIT distance="500" swimtime="00:07:56.27" />
                    <SPLIT distance="550" swimtime="00:08:45.09" />
                    <SPLIT distance="600" swimtime="00:09:35.15" />
                    <SPLIT distance="650" swimtime="00:10:23.06" />
                    <SPLIT distance="700" swimtime="00:11:12.48" />
                    <SPLIT distance="750" swimtime="00:12:00.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="334" swimtime="00:00:34.18" resultid="6662" heatid="10685" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1175" points="267" swimtime="00:03:15.69" resultid="6663" heatid="10716" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.05" />
                    <SPLIT distance="100" swimtime="00:01:33.65" />
                    <SPLIT distance="150" swimtime="00:02:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="265" swimtime="00:00:42.08" resultid="6664" heatid="10737" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="1287" points="305" swimtime="00:01:17.31" resultid="6665" heatid="10769" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="259" swimtime="00:00:38.29" resultid="6666" heatid="10822" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1467" points="273" swimtime="00:02:54.05" resultid="6667" heatid="10854" lane="1" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:24.84" />
                    <SPLIT distance="150" swimtime="00:02:11.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" status="DNS" swimtime="00:00:00.00" resultid="6668" heatid="10883" lane="5" entrytime="00:01:30.00" />
                <RESULT eventid="1674" status="DNS" swimtime="00:00:00.00" resultid="6669" heatid="10933" lane="7" entrytime="00:06:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-22" firstname="Alicja" gender="F" lastname="Romańska" nation="POL" athleteid="4211">
              <RESULTS>
                <RESULT eventid="1175" points="122" swimtime="00:04:13.73" resultid="6654" heatid="10713" lane="7" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.65" />
                    <SPLIT distance="100" swimtime="00:02:11.77" />
                    <SPLIT distance="150" swimtime="00:03:19.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="146" swimtime="00:04:23.84" resultid="6655" heatid="10752" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.04" />
                    <SPLIT distance="100" swimtime="00:02:11.91" />
                    <SPLIT distance="150" swimtime="00:03:19.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="58" swimtime="00:01:03.08" resultid="6656" heatid="10820" lane="6" entrytime="00:01:00.00" />
                <RESULT eventid="1467" points="128" swimtime="00:03:43.70" resultid="6657" heatid="10853" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.23" />
                    <SPLIT distance="100" swimtime="00:01:52.18" />
                    <SPLIT distance="150" swimtime="00:02:50.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="4172">
              <RESULTS>
                <RESULT eventid="1144" points="173" swimtime="00:00:42.57" resultid="6622" heatid="10681" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1175" points="37" swimtime="00:06:17.04" resultid="6623" heatid="10712" lane="4" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.76" />
                    <SPLIT distance="100" swimtime="00:03:14.34" />
                    <SPLIT distance="150" swimtime="00:04:56.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="62" swimtime="00:05:50.69" resultid="6624" heatid="10753" lane="0" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.58" />
                    <SPLIT distance="100" swimtime="00:02:48.99" />
                    <SPLIT distance="150" swimtime="00:04:22.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="45" swimtime="00:02:25.94" resultid="6625" heatid="10765" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="71" swimtime="00:02:35.30" resultid="6626" heatid="10803" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="22" swimtime="00:01:26.64" resultid="6627" heatid="10820" lane="7" entrytime="00:01:15.00" />
                <RESULT eventid="1562" points="25" swimtime="00:03:07.51" resultid="6628" heatid="10882" lane="3" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="81" swimtime="00:01:08.02" resultid="6629" heatid="10906" lane="0" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-03" firstname="Marcin" gender="M" lastname="Wyżga" nation="POL" athleteid="4207">
              <RESULTS>
                <RESULT eventid="1160" points="389" swimtime="00:00:28.64" resultid="6651" heatid="10704" lane="7" entrytime="00:00:28.50" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="6652" heatid="10782" lane="9" entrytime="00:01:04.50" />
                <RESULT eventid="1422" points="378" swimtime="00:00:31.01" resultid="6653" heatid="10833" lane="6" entrytime="00:00:30.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="4196">
              <RESULTS>
                <RESULT eventid="1098" points="85" swimtime="00:17:06.12" resultid="6642" heatid="10669" lane="8" entrytime="00:28:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.22" />
                    <SPLIT distance="100" swimtime="00:02:00.46" />
                    <SPLIT distance="150" swimtime="00:03:08.66" />
                    <SPLIT distance="200" swimtime="00:04:12.83" />
                    <SPLIT distance="250" swimtime="00:05:19.52" />
                    <SPLIT distance="300" swimtime="00:06:25.78" />
                    <SPLIT distance="350" swimtime="00:07:33.19" />
                    <SPLIT distance="400" swimtime="00:08:37.52" />
                    <SPLIT distance="450" swimtime="00:09:43.99" />
                    <SPLIT distance="500" swimtime="00:10:47.75" />
                    <SPLIT distance="550" swimtime="00:11:53.75" />
                    <SPLIT distance="600" swimtime="00:12:58.09" />
                    <SPLIT distance="650" swimtime="00:14:03.64" />
                    <SPLIT distance="700" swimtime="00:15:06.28" />
                    <SPLIT distance="750" swimtime="00:16:07.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="105" swimtime="00:00:44.28" resultid="6643" heatid="10691" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1302" points="96" swimtime="00:01:42.11" resultid="6644" heatid="10773" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="74" swimtime="00:04:02.63" resultid="6645" heatid="10857" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.44" />
                    <SPLIT distance="100" swimtime="00:01:52.98" />
                    <SPLIT distance="150" swimtime="00:02:57.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="71" swimtime="00:01:03.59" resultid="6646" heatid="10913" lane="1" entrytime="00:01:05.00" />
                <RESULT eventid="1695" points="79" swimtime="00:08:32.74" resultid="6647" heatid="10936" lane="7" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.12" />
                    <SPLIT distance="100" swimtime="00:02:00.63" />
                    <SPLIT distance="150" swimtime="00:03:08.60" />
                    <SPLIT distance="200" swimtime="00:04:15.28" />
                    <SPLIT distance="250" swimtime="00:05:23.03" />
                    <SPLIT distance="300" swimtime="00:06:28.35" />
                    <SPLIT distance="350" swimtime="00:07:32.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="4162">
              <RESULTS>
                <RESULT eventid="1128" points="136" swimtime="00:28:10.63" resultid="6613" heatid="10675" lane="5" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.11" />
                    <SPLIT distance="100" swimtime="00:01:48.76" />
                    <SPLIT distance="150" swimtime="00:02:45.61" />
                    <SPLIT distance="200" swimtime="00:03:42.96" />
                    <SPLIT distance="250" swimtime="00:04:40.42" />
                    <SPLIT distance="300" swimtime="00:05:37.79" />
                    <SPLIT distance="350" swimtime="00:06:34.88" />
                    <SPLIT distance="400" swimtime="00:07:32.24" />
                    <SPLIT distance="450" swimtime="00:08:29.19" />
                    <SPLIT distance="500" swimtime="00:09:25.63" />
                    <SPLIT distance="550" swimtime="00:10:21.07" />
                    <SPLIT distance="600" swimtime="00:11:17.28" />
                    <SPLIT distance="650" swimtime="00:12:13.35" />
                    <SPLIT distance="700" swimtime="00:13:09.81" />
                    <SPLIT distance="750" swimtime="00:14:06.38" />
                    <SPLIT distance="800" swimtime="00:15:02.13" />
                    <SPLIT distance="850" swimtime="00:15:57.33" />
                    <SPLIT distance="900" swimtime="00:16:53.95" />
                    <SPLIT distance="950" swimtime="00:17:49.89" />
                    <SPLIT distance="1000" swimtime="00:18:46.85" />
                    <SPLIT distance="1050" swimtime="00:19:44.12" />
                    <SPLIT distance="1100" swimtime="00:20:41.29" />
                    <SPLIT distance="1150" swimtime="00:21:38.73" />
                    <SPLIT distance="1200" swimtime="00:22:36.25" />
                    <SPLIT distance="1250" swimtime="00:23:33.35" />
                    <SPLIT distance="1300" swimtime="00:24:29.92" />
                    <SPLIT distance="1350" swimtime="00:25:27.38" />
                    <SPLIT distance="1400" swimtime="00:26:24.03" />
                    <SPLIT distance="1450" swimtime="00:27:20.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="196" swimtime="00:00:35.99" resultid="6614" heatid="10696" lane="6" entrytime="00:00:34.50" />
                <RESULT eventid="1190" points="113" swimtime="00:03:55.34" resultid="6615" heatid="10720" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.46" />
                    <SPLIT distance="100" swimtime="00:01:58.37" />
                    <SPLIT distance="150" swimtime="00:03:07.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="214" swimtime="00:01:18.37" resultid="6616" heatid="10777" lane="1" entrytime="00:01:16.00" />
                <RESULT eventid="1332" points="62" swimtime="00:04:40.25" resultid="6617" heatid="10792" lane="2" entrytime="00:04:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.23" />
                    <SPLIT distance="100" swimtime="00:02:13.28" />
                    <SPLIT distance="150" swimtime="00:03:23.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="157" swimtime="00:03:08.68" resultid="6618" heatid="10858" lane="6" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:01:29.45" />
                    <SPLIT distance="150" swimtime="00:02:20.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="97" swimtime="00:08:50.53" resultid="6619" heatid="10877" lane="8" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.62" />
                    <SPLIT distance="100" swimtime="00:02:05.81" />
                    <SPLIT distance="150" swimtime="00:03:18.63" />
                    <SPLIT distance="200" swimtime="00:04:31.59" />
                    <SPLIT distance="250" swimtime="00:05:43.08" />
                    <SPLIT distance="300" swimtime="00:06:57.30" />
                    <SPLIT distance="350" swimtime="00:07:55.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="79" swimtime="00:01:55.79" resultid="6620" heatid="10886" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="145" swimtime="00:06:58.43" resultid="6621" heatid="10937" lane="3" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                    <SPLIT distance="100" swimtime="00:01:45.26" />
                    <SPLIT distance="150" swimtime="00:02:40.96" />
                    <SPLIT distance="200" swimtime="00:03:36.82" />
                    <SPLIT distance="250" swimtime="00:04:30.36" />
                    <SPLIT distance="300" swimtime="00:05:23.47" />
                    <SPLIT distance="350" swimtime="00:06:12.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="4252">
              <RESULTS>
                <RESULT eventid="1160" points="326" swimtime="00:00:30.37" resultid="6689" heatid="10699" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1242" points="283" swimtime="00:00:36.59" resultid="6690" heatid="10747" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="6691" heatid="10779" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1422" points="379" swimtime="00:00:30.99" resultid="6692" heatid="10832" lane="9" entrytime="00:00:32.50" />
                <RESULT eventid="1452" points="266" swimtime="00:01:20.61" resultid="6693" heatid="10847" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="298" swimtime="00:01:14.53" resultid="6694" heatid="10888" lane="6" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="341" swimtime="00:00:37.81" resultid="6695" heatid="10919" lane="5" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="4242">
              <RESULTS>
                <RESULT eventid="1059" points="148" swimtime="00:15:14.85" resultid="6680" heatid="10666" lane="6" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                    <SPLIT distance="100" swimtime="00:01:41.02" />
                    <SPLIT distance="150" swimtime="00:02:41.36" />
                    <SPLIT distance="200" swimtime="00:03:38.67" />
                    <SPLIT distance="250" swimtime="00:04:37.57" />
                    <SPLIT distance="300" swimtime="00:05:34.86" />
                    <SPLIT distance="350" swimtime="00:06:32.52" />
                    <SPLIT distance="400" swimtime="00:07:30.54" />
                    <SPLIT distance="450" swimtime="00:08:29.19" />
                    <SPLIT distance="500" swimtime="00:09:27.25" />
                    <SPLIT distance="550" swimtime="00:10:24.83" />
                    <SPLIT distance="600" swimtime="00:11:22.23" />
                    <SPLIT distance="650" swimtime="00:12:08.76" />
                    <SPLIT distance="700" swimtime="00:13:19.01" />
                    <SPLIT distance="750" swimtime="00:14:18.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="245" swimtime="00:00:37.88" resultid="6681" heatid="10680" lane="4" />
                <RESULT eventid="1175" points="156" swimtime="00:03:54.20" resultid="6682" heatid="10714" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.30" />
                    <SPLIT distance="100" swimtime="00:01:52.51" />
                    <SPLIT distance="150" swimtime="00:03:00.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="203" swimtime="00:00:46.01" resultid="6683" heatid="10734" lane="0" />
                <RESULT eventid="1317" points="115" swimtime="00:04:10.29" resultid="6684" heatid="10789" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.37" />
                    <SPLIT distance="100" swimtime="00:01:58.95" />
                    <SPLIT distance="150" swimtime="00:03:05.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="156" swimtime="00:00:45.33" resultid="6685" heatid="10820" lane="8" />
                <RESULT eventid="1525" points="144" swimtime="00:08:27.60" resultid="6686" heatid="10873" lane="7" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.52" />
                    <SPLIT distance="100" swimtime="00:02:06.01" />
                    <SPLIT distance="150" swimtime="00:03:08.69" />
                    <SPLIT distance="200" swimtime="00:04:17.15" />
                    <SPLIT distance="250" swimtime="00:05:25.82" />
                    <SPLIT distance="300" swimtime="00:06:36.90" />
                    <SPLIT distance="350" swimtime="00:07:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="116" swimtime="00:01:53.64" resultid="6687" heatid="10882" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="136" swimtime="00:07:38.86" resultid="6688" heatid="10932" lane="1" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.65" />
                    <SPLIT distance="250" swimtime="00:04:42.91" />
                    <SPLIT distance="300" swimtime="00:05:42.21" />
                    <SPLIT distance="350" swimtime="00:06:41.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-09-18" firstname="Izabela" gender="F" lastname="Frączek" nation="POL" athleteid="4230">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat E 45-49  lat" eventid="1144" points="529" swimtime="00:00:29.33" resultid="6670" heatid="10688" lane="9" entrytime="00:00:29.60" />
                <RESULT eventid="1287" points="499" swimtime="00:01:05.62" resultid="6671" heatid="10770" lane="4" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat E  45-49  lat" eventid="1407" points="429" swimtime="00:00:32.37" resultid="6672" heatid="10824" lane="8" entrytime="00:00:32.95" />
                <RESULT eventid="1562" points="382" swimtime="00:01:16.45" resultid="6673" heatid="10884" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-21" firstname="Adam" gender="M" lastname="Pycia" nation="POL" athleteid="4181">
              <RESULTS>
                <RESULT eventid="1160" points="257" swimtime="00:00:32.86" resultid="6630" heatid="10698" lane="5" entrytime="00:00:31.50" />
                <RESULT eventid="1302" points="300" swimtime="00:01:10.02" resultid="6631" heatid="10779" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="251" swimtime="00:01:30.46" resultid="6632" heatid="10814" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="196" swimtime="00:00:38.61" resultid="6633" heatid="10828" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1638" points="294" swimtime="00:00:39.69" resultid="6634" heatid="10918" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="4235">
              <RESULTS>
                <RESULT eventid="1144" points="306" swimtime="00:00:35.20" resultid="6674" heatid="10683" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1175" points="223" swimtime="00:03:27.88" resultid="6675" heatid="10714" lane="0" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.55" />
                    <SPLIT distance="100" swimtime="00:01:42.80" />
                    <SPLIT distance="150" swimtime="00:02:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="236" swimtime="00:00:43.73" resultid="6676" heatid="10736" lane="9" entrytime="00:00:47.00" />
                <RESULT eventid="1407" points="242" swimtime="00:00:39.19" resultid="6677" heatid="10821" lane="6" entrytime="00:00:46.00" />
                <RESULT eventid="1437" points="217" swimtime="00:01:36.59" resultid="6678" heatid="10840" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="190" swimtime="00:03:35.55" resultid="6679" heatid="10895" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.02" />
                    <SPLIT distance="100" swimtime="00:01:49.66" />
                    <SPLIT distance="150" swimtime="00:02:47.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" name="Korona Kraków C" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="359" swimtime="00:02:11.45" resultid="6699" heatid="10801" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:13.23" />
                    <SPLIT distance="150" swimtime="00:01:43.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4252" number="1" />
                    <RELAYPOSITION athleteid="4158" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4216" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4207" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" name="Korona Kraków D" number="1">
              <RESULTS>
                <RESULT eventid="1518" points="319" swimtime="00:02:04.14" resultid="6703" heatid="10871" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:36.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4181" number="1" />
                    <RELAYPOSITION athleteid="4158" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4162" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4207" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" name="Korona Kraków E" number="2">
              <RESULTS>
                <RESULT eventid="1368" points="170" swimtime="00:02:48.53" resultid="6700" heatid="10800" lane="7" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.84" />
                    <SPLIT distance="100" swimtime="00:01:33.17" />
                    <SPLIT distance="150" swimtime="00:02:04.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4162" number="1" />
                    <RELAYPOSITION athleteid="4181" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4187" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4196" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F" name="Korona Kraków D" number="1">
              <RESULTS>
                <RESULT eventid="1347" points="386" swimtime="00:02:26.00" resultid="6701" heatid="10798" lane="6" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:01:20.25" />
                    <SPLIT distance="150" swimtime="00:01:57.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4220" number="1" />
                    <RELAYPOSITION athleteid="4151" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4203" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4230" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters w  kat D  200-239  lat" eventid="1497" points="426" swimtime="00:02:08.19" resultid="6702" heatid="10868" lane="2" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                    <SPLIT distance="100" swimtime="00:01:03.39" />
                    <SPLIT distance="150" swimtime="00:01:38.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4230" number="1" />
                    <RELAYPOSITION athleteid="4203" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4220" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4151" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="Korona Kraków C" number="1">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  w  kat C  160-199  lat" eventid="1205" swimtime="00:01:53.30" resultid="6696" heatid="10733" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="100" swimtime="00:00:58.23" />
                    <SPLIT distance="150" swimtime="00:01:26.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4151" number="1" />
                    <RELAYPOSITION athleteid="4207" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4230" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4216" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1653" swimtime="00:02:14.12" resultid="6697" heatid="10929" lane="0" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:01:14.80" />
                    <SPLIT distance="150" swimtime="00:01:45.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4151" number="1" />
                    <RELAYPOSITION athleteid="4158" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4207" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4230" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" name="Korona Kraków D" number="2">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:11.45" resultid="6698" heatid="10732" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:02.04" />
                    <SPLIT distance="150" swimtime="00:01:36.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4181" number="1" />
                    <RELAYPOSITION athleteid="4187" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4220" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4203" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" name="Korona Kraków E" number="2">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:46.37" resultid="6704" heatid="10928" lane="8" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.50" />
                    <SPLIT distance="100" swimtime="00:01:24.04" />
                    <SPLIT distance="150" swimtime="00:02:01.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4242" number="1" />
                    <RELAYPOSITION athleteid="4252" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4203" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4196" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KPPOL" nation="POL" region="14" clubid="5615" name="KPMG Polska">
          <CONTACT name="s" />
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Piotr" gender="M" lastname="Kotynia" nation="POL" athleteid="5629">
              <RESULTS>
                <RESULT eventid="1160" points="368" swimtime="00:00:29.16" resultid="7136" heatid="10709" lane="0" entrytime="00:00:26.30" />
                <RESULT eventid="1272" points="317" swimtime="00:03:06.15" resultid="7137" heatid="10764" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:23.13" />
                    <SPLIT distance="150" swimtime="00:02:13.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="335" swimtime="00:01:22.18" resultid="7138" heatid="10819" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="362" swimtime="00:00:31.46" resultid="7139" heatid="10836" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="1638" points="426" swimtime="00:00:35.10" resultid="7140" heatid="10926" lane="1" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Patryk" gender="M" lastname="Bednarz" nation="POL" athleteid="5623">
              <RESULTS>
                <RESULT eventid="1160" points="316" swimtime="00:00:30.68" resultid="7131" heatid="10700" lane="7" entrytime="00:00:30.16" />
                <RESULT eventid="1302" points="320" swimtime="00:01:08.57" resultid="7132" heatid="10780" lane="9" entrytime="00:01:08.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="312" swimtime="00:00:33.04" resultid="7133" heatid="10829" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1482" points="289" swimtime="00:02:34.19" resultid="7134" heatid="10861" lane="9" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                    <SPLIT distance="150" swimtime="00:01:55.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="214" swimtime="00:01:23.27" resultid="7135" heatid="10888" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Adam" gender="M" lastname="Heromiński" nation="POL" athleteid="5635">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="7141" heatid="10691" lane="2" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NERZI" nation="SVK" clubid="10657" name="KPS Nereus Zilina">
          <ATHLETES>
            <ATHLETE birthdate="1960-01-01" firstname="Rastislav" gender="M" lastname="Pavlik" nation="POL" athleteid="7310">
              <RESULTS>
                <RESULT eventid="1160" points="416" swimtime="00:00:27.99" resultid="9916" heatid="10705" lane="6" entrytime="00:00:27.86" />
                <RESULT eventid="1242" points="394" swimtime="00:00:32.77" resultid="9917" heatid="10749" lane="7" entrytime="00:00:32.23" />
                <RESULT eventid="1302" points="399" swimtime="00:01:03.70" resultid="9918" heatid="10782" lane="4" entrytime="00:01:03.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="365" swimtime="00:01:12.55" resultid="9919" heatid="10849" lane="9" entrytime="00:01:10.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="329" swimtime="00:02:42.12" resultid="9920" heatid="10903" lane="6" entrytime="00:02:38.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:19.13" />
                    <SPLIT distance="150" swimtime="00:02:01.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="343" swimtime="00:00:37.72" resultid="9921" heatid="10923" lane="1" entrytime="00:00:35.23" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" region="EXOBO" clubid="2895" name="Ks Extreme Team Oborniki">
          <CONTACT city="OBORNIKI" email="JANWOL@POCZTA.ONET.PL" name="WOLNIEWICZ JANUSZ" phone="791064667" state="WIE" street="CZARNKOWSKA 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="2896">
              <RESULTS>
                <RESULT eventid="1128" points="99" swimtime="00:31:22.20" resultid="7550" heatid="10675" lane="7" entrytime="00:28:53.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.96" />
                    <SPLIT distance="100" swimtime="00:01:49.20" />
                    <SPLIT distance="150" swimtime="00:02:49.33" />
                    <SPLIT distance="200" swimtime="00:03:49.81" />
                    <SPLIT distance="250" swimtime="00:04:51.01" />
                    <SPLIT distance="350" swimtime="00:05:13.18" />
                    <SPLIT distance="400" swimtime="00:05:53.08" />
                    <SPLIT distance="450" swimtime="00:06:55.49" />
                    <SPLIT distance="500" swimtime="00:07:58.68" />
                    <SPLIT distance="550" swimtime="00:09:01.25" />
                    <SPLIT distance="600" swimtime="00:10:04.74" />
                    <SPLIT distance="650" swimtime="00:11:07.86" />
                    <SPLIT distance="700" swimtime="00:12:11.04" />
                    <SPLIT distance="750" swimtime="00:13:15.71" />
                    <SPLIT distance="850" swimtime="00:13:48.16" />
                    <SPLIT distance="900" swimtime="00:14:20.70" />
                    <SPLIT distance="950" swimtime="00:15:25.27" />
                    <SPLIT distance="1000" swimtime="00:16:29.16" />
                    <SPLIT distance="1050" swimtime="00:17:33.01" />
                    <SPLIT distance="1100" swimtime="00:18:37.47" />
                    <SPLIT distance="1150" swimtime="00:19:41.18" />
                    <SPLIT distance="1200" swimtime="00:20:45.50" />
                    <SPLIT distance="1250" swimtime="00:21:49.41" />
                    <SPLIT distance="1300" swimtime="00:22:53.04" />
                    <SPLIT distance="1350" swimtime="00:23:55.74" />
                    <SPLIT distance="1400" swimtime="00:24:58.86" />
                    <SPLIT distance="1450" swimtime="00:26:03.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="7551" heatid="10694" lane="9" entrytime="00:00:36.15" entrycourse="SCM" />
                <RESULT eventid="1302" points="150" swimtime="00:01:28.23" resultid="7552" heatid="10775" lane="1" entrytime="00:01:23.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="111" swimtime="00:03:31.77" resultid="7553" heatid="10857" lane="4" entrytime="00:03:18.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="100" swimtime="00:01:39.13" />
                    <SPLIT distance="150" swimtime="00:02:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="100" swimtime="00:07:52.67" resultid="7554" heatid="10937" lane="9" entrytime="00:07:15.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.68" />
                    <SPLIT distance="100" swimtime="00:01:49.41" />
                    <SPLIT distance="150" swimtime="00:02:50.09" />
                    <SPLIT distance="200" swimtime="00:03:52.31" />
                    <SPLIT distance="250" swimtime="00:04:53.90" />
                    <SPLIT distance="300" swimtime="00:05:54.73" />
                    <SPLIT distance="350" swimtime="00:06:56.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GORAD" nation="POL" region="SLA" clubid="3403" name="Ks Górnik Radlin 00211">
          <CONTACT name="CYMERMAN IWONA" />
          <ATHLETES>
            <ATHLETE birthdate="1985-11-07" firstname="Iwona" gender="F" lastname="Cymerman" nation="POL" athleteid="3409">
              <RESULTS>
                <RESULT eventid="1287" points="472" swimtime="00:01:06.85" resultid="7935" heatid="10771" lane="9" entrytime="00:01:06.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="421" swimtime="00:00:32.59" resultid="7936" heatid="10824" lane="1" entrytime="00:00:32.86" />
                <RESULT eventid="1467" points="369" swimtime="00:02:37.50" resultid="7937" heatid="10855" lane="0" entrytime="00:02:33.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:13.24" />
                    <SPLIT distance="150" swimtime="00:01:55.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="435" swimtime="00:00:38.89" resultid="7938" heatid="10910" lane="5" entrytime="00:00:39.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MYDAB" nation="POL" region="SLA" clubid="3620" name="KS Mydlice Dąbrowa Górnicza">
          <CONTACT name="s" />
          <ATHLETES>
            <ATHLETE birthdate="1996-01-01" firstname="Mateusz" gender="M" lastname="Burzawa" nation="POL" athleteid="3621">
              <RESULTS>
                <RESULT eventid="1098" points="407" swimtime="00:10:09.60" resultid="3622" heatid="10668" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                    <SPLIT distance="150" swimtime="00:01:46.19" />
                    <SPLIT distance="200" swimtime="00:02:24.38" />
                    <SPLIT distance="250" swimtime="00:03:03.04" />
                    <SPLIT distance="300" swimtime="00:03:41.62" />
                    <SPLIT distance="350" swimtime="00:04:20.46" />
                    <SPLIT distance="400" swimtime="00:04:59.55" />
                    <SPLIT distance="450" swimtime="00:05:39.08" />
                    <SPLIT distance="500" swimtime="00:06:18.94" />
                    <SPLIT distance="550" swimtime="00:06:58.77" />
                    <SPLIT distance="600" swimtime="00:07:38.13" />
                    <SPLIT distance="650" swimtime="00:08:17.12" />
                    <SPLIT distance="700" swimtime="00:08:56.04" />
                    <SPLIT distance="750" swimtime="00:09:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="489" swimtime="00:02:24.61" resultid="3623" heatid="10729" lane="3" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                    <SPLIT distance="100" swimtime="00:01:08.94" />
                    <SPLIT distance="150" swimtime="00:01:51.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="3624" heatid="10750" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1272" points="422" swimtime="00:02:49.32" resultid="3625" heatid="10764" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                    <SPLIT distance="100" swimtime="00:01:20.95" />
                    <SPLIT distance="150" swimtime="00:02:05.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="3626" heatid="10818" lane="4" entrytime="00:01:13.00" />
                <RESULT eventid="1452" status="DNS" swimtime="00:00:00.00" resultid="3627" heatid="10849" lane="2" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="DOL" clubid="5218" name="Ks Rekin Świebodzice">
          <CONTACT city="Świebodzice" email="winiar182@wp.pl" internet="www.klubrekin.pl" name="WINIARCZYK Krzysztof" phone="606626274" state="DOL" street="Mieszka Starego 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1982-11-09" firstname="Karol" gender="M" lastname="Żemier" nation="POL" athleteid="9879">
              <RESULTS>
                <RESULT eventid="1160" points="501" swimtime="00:00:26.32" resultid="9880" heatid="10689" lane="8" />
                <RESULT eventid="1190" points="464" swimtime="00:02:27.18" resultid="9881" heatid="10730" lane="9" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:51.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="524" swimtime="00:00:29.81" resultid="9882" heatid="10751" lane="2" entrytime="00:00:28.60" />
                <RESULT eventid="1332" points="413" swimtime="00:02:29.67" resultid="9883" heatid="10796" lane="6" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:10.16" />
                    <SPLIT distance="150" swimtime="00:01:49.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="540" swimtime="00:00:27.53" resultid="9884" heatid="10826" lane="8" />
                <RESULT eventid="1452" points="502" swimtime="00:01:05.20" resultid="9885" heatid="10850" lane="2" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="517" swimtime="00:01:02.06" resultid="9886" heatid="10885" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="429" swimtime="00:02:28.36" resultid="9887" heatid="10898" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:10.54" />
                    <SPLIT distance="150" swimtime="00:01:50.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-18" firstname="Marek" gender="M" lastname="Stuczyński" nation="POL" athleteid="9874">
              <RESULTS>
                <RESULT eventid="1160" points="513" swimtime="00:00:26.12" resultid="9875" heatid="10710" lane="9" entrytime="00:00:25.50" entrycourse="SCM" />
                <RESULT eventid="1302" points="497" swimtime="00:00:59.22" resultid="9876" heatid="10787" lane="0" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="430" swimtime="00:01:15.67" resultid="9877" heatid="10819" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="574" swimtime="00:00:31.78" resultid="9878" heatid="10926" lane="8" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-21" firstname="Alfred" gender="M" lastname="Żemier" nation="POL" athleteid="9888">
              <RESULTS>
                <RESULT eventid="1160" points="487" swimtime="00:00:26.57" resultid="9889" heatid="10690" lane="7" />
                <RESULT eventid="1190" points="343" swimtime="00:02:42.85" resultid="9890" heatid="10727" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:02:04.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="424" swimtime="00:00:31.98" resultid="9891" heatid="10750" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1302" points="468" swimtime="00:01:00.39" resultid="9892" heatid="10784" lane="7" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="475" swimtime="00:00:28.74" resultid="9893" heatid="10826" lane="1" />
                <RESULT eventid="1452" points="379" swimtime="00:01:11.59" resultid="9894" heatid="10850" lane="8" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="334" swimtime="00:02:41.21" resultid="9895" heatid="10899" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:19.43" />
                    <SPLIT distance="150" swimtime="00:02:01.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-12-12" firstname="Karolina" gender="F" lastname="Jahnz" nation="POL" athleteid="9856">
              <RESULTS>
                <RESULT eventid="1113" points="322" swimtime="00:22:29.04" resultid="9857" heatid="10674" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="150" swimtime="00:02:06.07" />
                    <SPLIT distance="200" swimtime="00:02:51.64" />
                    <SPLIT distance="250" swimtime="00:03:37.02" />
                    <SPLIT distance="300" swimtime="00:04:22.43" />
                    <SPLIT distance="350" swimtime="00:05:07.80" />
                    <SPLIT distance="400" swimtime="00:05:53.38" />
                    <SPLIT distance="450" swimtime="00:06:38.39" />
                    <SPLIT distance="500" swimtime="00:07:23.81" />
                    <SPLIT distance="550" swimtime="00:08:09.31" />
                    <SPLIT distance="600" swimtime="00:08:54.58" />
                    <SPLIT distance="650" swimtime="00:09:40.18" />
                    <SPLIT distance="700" swimtime="00:10:25.36" />
                    <SPLIT distance="750" swimtime="00:11:10.69" />
                    <SPLIT distance="800" swimtime="00:11:56.22" />
                    <SPLIT distance="850" swimtime="00:12:41.56" />
                    <SPLIT distance="900" swimtime="00:13:27.17" />
                    <SPLIT distance="950" swimtime="00:14:12.41" />
                    <SPLIT distance="1000" swimtime="00:14:57.93" />
                    <SPLIT distance="1050" swimtime="00:15:42.94" />
                    <SPLIT distance="1100" swimtime="00:16:28.40" />
                    <SPLIT distance="1150" swimtime="00:17:14.30" />
                    <SPLIT distance="1200" swimtime="00:17:59.88" />
                    <SPLIT distance="1250" swimtime="00:18:45.26" />
                    <SPLIT distance="1300" swimtime="00:19:30.58" />
                    <SPLIT distance="1350" swimtime="00:20:16.45" />
                    <SPLIT distance="1400" swimtime="00:21:01.12" />
                    <SPLIT distance="1450" swimtime="00:21:45.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="345" swimtime="00:02:59.78" resultid="9858" heatid="10712" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="100" swimtime="00:01:26.68" />
                    <SPLIT distance="150" swimtime="00:02:18.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="319" swimtime="00:03:23.49" resultid="9859" heatid="10752" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                    <SPLIT distance="100" swimtime="00:01:38.64" />
                    <SPLIT distance="150" swimtime="00:02:31.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1317" points="240" swimtime="00:03:15.90" resultid="9860" heatid="10790" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:31.47" />
                    <SPLIT distance="150" swimtime="00:02:23.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="357" swimtime="00:02:39.20" resultid="9861" heatid="10851" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:15.93" />
                    <SPLIT distance="150" swimtime="00:01:58.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="357" swimtime="00:06:15.45" resultid="9862" heatid="10874" lane="5" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:31.31" />
                    <SPLIT distance="150" swimtime="00:02:20.87" />
                    <SPLIT distance="200" swimtime="00:03:08.29" />
                    <SPLIT distance="250" swimtime="00:04:00.89" />
                    <SPLIT distance="300" swimtime="00:04:53.34" />
                    <SPLIT distance="350" swimtime="00:05:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="325" swimtime="00:03:00.34" resultid="9863" heatid="10893" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                    <SPLIT distance="100" swimtime="00:01:26.79" />
                    <SPLIT distance="150" swimtime="00:02:14.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="364" swimtime="00:05:30.94" resultid="9864" heatid="10933" lane="2" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                    <SPLIT distance="100" swimtime="00:01:17.67" />
                    <SPLIT distance="150" swimtime="00:02:00.28" />
                    <SPLIT distance="200" swimtime="00:02:43.29" />
                    <SPLIT distance="250" swimtime="00:03:25.96" />
                    <SPLIT distance="300" swimtime="00:04:09.08" />
                    <SPLIT distance="350" swimtime="00:04:51.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-13" firstname="Magdalena" gender="F" lastname="Stachowska" nation="POL" athleteid="9865">
              <RESULTS>
                <RESULT eventid="1059" points="199" swimtime="00:13:49.94" resultid="9866" heatid="10665" lane="5" />
                <RESULT eventid="1144" points="380" swimtime="00:00:32.74" resultid="9867" heatid="10687" lane="0" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1175" points="223" swimtime="00:03:27.77" resultid="9868" heatid="10712" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="100" swimtime="00:01:41.04" />
                    <SPLIT distance="150" swimtime="00:02:40.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="239" swimtime="00:03:43.92" resultid="9869" heatid="10752" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.16" />
                    <SPLIT distance="100" swimtime="00:01:49.85" />
                    <SPLIT distance="150" swimtime="00:02:48.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="302" swimtime="00:01:17.58" resultid="9870" heatid="10770" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="281" swimtime="00:01:38.17" resultid="9871" heatid="10807" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="214" swimtime="00:03:08.82" resultid="9872" heatid="10851" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="100" swimtime="00:01:26.67" />
                    <SPLIT distance="150" swimtime="00:02:18.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="335" swimtime="00:00:42.43" resultid="9873" heatid="10909" lane="6" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-22" firstname="Aleksandra" gender="F" lastname="Hebel" nation="POL" athleteid="9848">
              <RESULTS>
                <RESULT eventid="1144" points="375" swimtime="00:00:32.89" resultid="9849" heatid="10686" lane="8" entrytime="00:00:33.50" entrycourse="SCM" />
                <RESULT eventid="1257" points="227" swimtime="00:03:47.71" resultid="9850" heatid="10752" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.05" />
                    <SPLIT distance="100" swimtime="00:01:49.58" />
                    <SPLIT distance="150" swimtime="00:02:48.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="328" swimtime="00:01:15.47" resultid="9851" heatid="10769" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="225" swimtime="00:01:45.74" resultid="9852" heatid="10806" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="277" swimtime="00:02:53.17" resultid="9853" heatid="10853" lane="6" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:22.70" />
                    <SPLIT distance="150" swimtime="00:02:09.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="259" swimtime="00:03:14.59" resultid="9854" heatid="10895" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.70" />
                    <SPLIT distance="100" swimtime="00:01:35.16" />
                    <SPLIT distance="150" swimtime="00:02:25.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="213" swimtime="00:00:49.33" resultid="9855" heatid="10908" lane="9" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-20" firstname="Veronica" gender="F" lastname="Campbell-Żemier" nation="POL" athleteid="9843">
              <RESULTS>
                <RESULT eventid="1144" points="504" swimtime="00:00:29.80" resultid="9844" heatid="10686" lane="3" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1287" points="501" swimtime="00:01:05.53" resultid="9845" heatid="10768" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="411" swimtime="00:01:26.53" resultid="9846" heatid="10807" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="431" swimtime="00:00:39.02" resultid="9847" heatid="10911" lane="7" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-16" firstname="Filip" gender="M" lastname="Żemier" nation="POL" athleteid="9896">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="9897" heatid="10708" lane="1" entrytime="00:00:26.90" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="9898" heatid="10782" lane="3" entrytime="00:01:03.50" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="9899" heatid="10835" lane="0" entrytime="00:00:29.90" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="9900" heatid="10891" lane="8" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" name="Rekin Świebodzice" number="1">
              <RESULTS>
                <RESULT eventid="1518" status="DNS" swimtime="00:00:00.00" resultid="9901" heatid="10869" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9843" number="1" />
                    <RELAYPOSITION athleteid="9874" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9848" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9879" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" name="Rekin Świebodzice" number="1">
              <RESULTS>
                <RESULT eventid="1347" points="334" swimtime="00:02:33.10" resultid="9903" heatid="10798" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:24.76" />
                    <SPLIT distance="150" swimtime="00:02:03.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9865" number="1" />
                    <RELAYPOSITION athleteid="9843" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9856" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9848" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1497" points="433" swimtime="00:02:07.58" resultid="9904" heatid="10868" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:03.10" />
                    <SPLIT distance="150" swimtime="00:01:35.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9843" number="1" />
                    <RELAYPOSITION athleteid="9848" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9856" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9865" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="Rekin Świebodzice" number="1">
              <RESULTS>
                <RESULT eventid="1653" status="DNS" swimtime="00:00:00.00" resultid="9902" heatid="10929" lane="2" entrytime="00:02:08.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9879" number="1" />
                    <RELAYPOSITION athleteid="9874" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9865" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9843" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1205" swimtime="00:01:57.89" resultid="9905" heatid="10733" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                    <SPLIT distance="100" swimtime="00:00:59.11" />
                    <SPLIT distance="150" swimtime="00:01:31.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9874" number="1" />
                    <RELAYPOSITION athleteid="9848" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9856" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9896" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1653" status="DNS" swimtime="00:00:00.00" resultid="9906" heatid="10928" lane="2" entrytime="00:02:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9888" number="1" />
                    <RELAYPOSITION athleteid="9856" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9896" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9848" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1653" swimtime="00:02:08.23" resultid="9908" heatid="10929" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="100" swimtime="00:01:07.81" />
                    <SPLIT distance="150" swimtime="00:01:36.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9879" number="1" />
                    <RELAYPOSITION athleteid="9865" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9888" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9843" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" name="Rekin Świebodzice" number="2">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="9907" heatid="10733" lane="4" entrytime="00:01:50.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9874" number="1" />
                    <RELAYPOSITION athleteid="9888" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9896" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9879" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="15" clubid="9370" name="KU AZS UAM Poznań">
          <CONTACT city="Poznań" email="kukowalazs@gmail.com" name="Kowalik" phone="603965223" state="WLKP" street="Zagajnikowa 9" zip="61-602" />
          <ATHLETES>
            <ATHLETE birthdate="1981-12-27" firstname="Bartosz" gender="M" lastname="Jankowiak" nation="POL" athleteid="9371">
              <RESULTS>
                <RESULT eventid="1128" points="253" swimtime="00:22:56.09" resultid="9372" heatid="10678" lane="9" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:02:07.22" />
                    <SPLIT distance="200" swimtime="00:02:53.16" />
                    <SPLIT distance="250" swimtime="00:03:39.12" />
                    <SPLIT distance="300" swimtime="00:04:25.28" />
                    <SPLIT distance="350" swimtime="00:05:11.31" />
                    <SPLIT distance="400" swimtime="00:05:57.16" />
                    <SPLIT distance="450" swimtime="00:06:43.14" />
                    <SPLIT distance="500" swimtime="00:07:29.23" />
                    <SPLIT distance="550" swimtime="00:08:15.61" />
                    <SPLIT distance="600" swimtime="00:09:01.81" />
                    <SPLIT distance="650" swimtime="00:09:48.38" />
                    <SPLIT distance="700" swimtime="00:10:34.87" />
                    <SPLIT distance="750" swimtime="00:11:21.68" />
                    <SPLIT distance="800" swimtime="00:12:08.03" />
                    <SPLIT distance="850" swimtime="00:12:54.41" />
                    <SPLIT distance="900" swimtime="00:13:41.13" />
                    <SPLIT distance="950" swimtime="00:14:27.86" />
                    <SPLIT distance="1000" swimtime="00:15:14.64" />
                    <SPLIT distance="1050" swimtime="00:16:01.02" />
                    <SPLIT distance="1100" swimtime="00:16:48.16" />
                    <SPLIT distance="1150" swimtime="00:17:34.60" />
                    <SPLIT distance="1200" swimtime="00:18:21.20" />
                    <SPLIT distance="1250" swimtime="00:19:07.59" />
                    <SPLIT distance="1300" swimtime="00:19:54.12" />
                    <SPLIT distance="1350" swimtime="00:20:40.93" />
                    <SPLIT distance="1400" swimtime="00:21:27.47" />
                    <SPLIT distance="1450" swimtime="00:22:13.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UW" nation="POL" region="14" clubid="5637" name="KU AZS Uniwersytet Warszawski">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1993-01-01" firstname="Krzysztof" gender="M" lastname="Micorek" nation="POL" athleteid="5638">
              <RESULTS>
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="7146" heatid="10740" lane="5" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="7147" heatid="10772" lane="3" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="7148" heatid="10825" lane="3" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="7149" heatid="10885" lane="1" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="7150" heatid="10912" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LAFUR" nation="POL" region="MAZ" clubid="9376" name="Laguna Furmana">
          <CONTACT city="WARSZAWA" name="FURMAN PIOTR" phone="602655550" state="MAZ" street="PODLEŚNA 40/26" zip="01-673" />
          <ATHLETES>
            <ATHLETE birthdate="1961-03-18" firstname="Piotr" gender="M" lastname="Furman" nation="POL" athleteid="9377">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="9378" heatid="10703" lane="5" entrytime="00:00:28.99" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="9379" heatid="10830" lane="3" entrytime="00:00:33.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06614" nation="POL" region="14" clubid="4306" name="Legia Warszawa">
          <CONTACT email="janek@plywanielegia.pl" name="Peńsko" phone="600826305" />
          <ATHLETES>
            <ATHLETE birthdate="1981-10-24" firstname="Marcin" gender="M" lastname="wilczęga" nation="POL" athleteid="4347">
              <RESULTS>
                <RESULT eventid="1160" points="432" swimtime="00:00:27.65" resultid="6809" heatid="10689" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="4307">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Mężczyzn w  kat D  40-44  lata" eventid="1160" points="551" swimtime="00:00:25.50" resultid="6776" heatid="10689" lane="3" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn  w  kat D  40-44  lata" eventid="1242" points="615" swimtime="00:00:28.26" resultid="6777" heatid="10751" lane="7" entrytime="00:00:28.80" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn  w  kat D  40-44  lat" eventid="1422" points="614" swimtime="00:00:26.38" resultid="6778" heatid="10825" lane="4" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn w  kat D  40-44  lat" eventid="1452" points="581" swimtime="00:01:02.11" resultid="6779" heatid="10850" lane="3" entrytime="00:01:02.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1578" points="593" swimtime="00:00:59.27" resultid="6780" heatid="10892" lane="2" entrytime="00:00:59.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-07" firstname="Agnieszka" gender="F" lastname="Kaczmarek" nation="POL" athleteid="4313">
              <RESULTS>
                <RESULT eventid="1144" points="519" swimtime="00:00:29.52" resultid="6781" heatid="10685" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1175" points="488" swimtime="00:02:40.15" resultid="6782" heatid="10718" lane="7" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:15.57" />
                    <SPLIT distance="150" swimtime="00:02:00.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat B  30-34  lat" eventid="1226" points="527" swimtime="00:00:33.49" resultid="6783" heatid="10739" lane="7" entrytime="00:00:33.50" />
                <RESULT eventid="1407" status="DNS" swimtime="00:00:00.00" resultid="6784" heatid="10820" lane="1" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat B  30-34  lata" eventid="1437" points="511" swimtime="00:01:12.67" resultid="6785" heatid="10842" lane="6" entrytime="00:01:13.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" status="DNS" swimtime="00:00:00.00" resultid="6786" heatid="10882" lane="2" />
                <RESULT eventid="1623" points="436" swimtime="00:00:38.85" resultid="6787" heatid="10908" lane="7" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-12" firstname="Filip" gender="M" lastname="Rowiński" nation="POL" athleteid="4354">
              <RESULTS>
                <RESULT eventid="1160" points="519" swimtime="00:00:26.01" resultid="6813" heatid="10689" lane="9" />
                <RESULT eventid="1272" points="576" swimtime="00:02:32.65" resultid="6814" heatid="10764" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:12.79" />
                    <SPLIT distance="150" swimtime="00:01:53.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="573" swimtime="00:00:27.00" resultid="6815" heatid="10837" lane="8" entrytime="00:00:28.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1638" points="710" swimtime="00:00:29.61" resultid="6817" heatid="10926" lane="6" entrytime="00:00:29.70" />
                <RESULT eventid="1392" points="632" swimtime="00:01:06.57" resultid="9531" heatid="10819" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-21" firstname="Krzysztof" gender="M" lastname="Spyra" nation="POL" athleteid="4351">
              <RESULTS>
                <RESULT eventid="1160" points="434" swimtime="00:00:27.61" resultid="6811" heatid="10689" lane="7" />
                <RESULT eventid="1695" points="403" swimtime="00:04:57.71" resultid="6812" heatid="10935" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:08.82" />
                    <SPLIT distance="150" swimtime="00:01:46.14" />
                    <SPLIT distance="200" swimtime="00:02:23.77" />
                    <SPLIT distance="250" swimtime="00:03:01.82" />
                    <SPLIT distance="300" swimtime="00:03:40.55" />
                    <SPLIT distance="350" swimtime="00:04:19.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-13" firstname="Paweł" gender="M" lastname="Korzeniowski" nation="POL" athleteid="4333">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Mężczyzn w  kat B  30-34 lata" eventid="1160" points="707" swimtime="00:00:23.47" resultid="6798" heatid="10689" lane="4" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn w  kat B  30-34  lata" eventid="1302" points="782" swimtime="00:00:50.91" resultid="6799" heatid="10788" lane="4" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="4321">
              <RESULTS>
                <RESULT eventid="1160" points="237" swimtime="00:00:33.77" resultid="6788" heatid="10697" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1190" points="158" swimtime="00:03:30.56" resultid="6789" heatid="10721" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                    <SPLIT distance="100" swimtime="00:01:40.78" />
                    <SPLIT distance="150" swimtime="00:02:44.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="200" swimtime="00:00:41.05" resultid="6790" heatid="10744" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1332" points="85" swimtime="00:04:13.08" resultid="6791" heatid="10792" lane="3" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.46" />
                    <SPLIT distance="100" swimtime="00:02:01.53" />
                    <SPLIT distance="150" swimtime="00:03:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="163" swimtime="00:01:34.80" resultid="6792" heatid="10845" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="141" swimtime="00:07:47.91" resultid="6793" heatid="10877" lane="1" entrytime="00:07:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="150" swimtime="00:00:56.00" />
                    <SPLIT distance="200" swimtime="00:03:55.31" />
                    <SPLIT distance="250" swimtime="00:05:03.41" />
                    <SPLIT distance="300" swimtime="00:06:11.93" />
                    <SPLIT distance="350" swimtime="00:07:01.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="140" swimtime="00:03:35.28" resultid="6794" heatid="10900" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.08" />
                    <SPLIT distance="100" swimtime="00:01:46.25" />
                    <SPLIT distance="150" swimtime="00:02:41.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="188" swimtime="00:06:23.97" resultid="6795" heatid="10938" lane="1" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:29.31" />
                    <SPLIT distance="150" swimtime="00:02:18.50" />
                    <SPLIT distance="200" swimtime="00:03:08.89" />
                    <SPLIT distance="250" swimtime="00:04:00.70" />
                    <SPLIT distance="300" swimtime="00:04:50.69" />
                    <SPLIT distance="350" swimtime="00:05:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="177" swimtime="00:25:49.97" resultid="9803" heatid="10675" lane="2" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:29.81" />
                    <SPLIT distance="150" swimtime="00:02:19.29" />
                    <SPLIT distance="200" swimtime="00:03:11.00" />
                    <SPLIT distance="250" swimtime="00:04:02.80" />
                    <SPLIT distance="300" swimtime="00:04:55.74" />
                    <SPLIT distance="350" swimtime="00:05:48.40" />
                    <SPLIT distance="400" swimtime="00:06:41.59" />
                    <SPLIT distance="450" swimtime="00:07:35.63" />
                    <SPLIT distance="500" swimtime="00:08:28.94" />
                    <SPLIT distance="550" swimtime="00:09:22.78" />
                    <SPLIT distance="600" swimtime="00:10:15.70" />
                    <SPLIT distance="650" swimtime="00:11:07.85" />
                    <SPLIT distance="700" swimtime="00:12:00.36" />
                    <SPLIT distance="750" swimtime="00:12:52.55" />
                    <SPLIT distance="800" swimtime="00:13:44.71" />
                    <SPLIT distance="850" swimtime="00:14:37.06" />
                    <SPLIT distance="900" swimtime="00:15:30.20" />
                    <SPLIT distance="950" swimtime="00:16:23.27" />
                    <SPLIT distance="1000" swimtime="00:17:15.82" />
                    <SPLIT distance="1050" swimtime="00:18:08.03" />
                    <SPLIT distance="1100" swimtime="00:19:00.53" />
                    <SPLIT distance="1150" swimtime="00:19:52.59" />
                    <SPLIT distance="1200" swimtime="00:20:44.64" />
                    <SPLIT distance="1250" swimtime="00:21:36.45" />
                    <SPLIT distance="1300" swimtime="00:22:28.82" />
                    <SPLIT distance="1350" swimtime="00:23:21.56" />
                    <SPLIT distance="1400" swimtime="00:24:13.43" />
                    <SPLIT distance="1450" swimtime="00:25:03.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-16" firstname="Jacek" gender="M" lastname="Kaczyński" nation="POL" athleteid="4330">
              <RESULTS>
                <RESULT eventid="1160" points="656" swimtime="00:00:24.06" resultid="6796" heatid="10689" lane="5" />
                <RESULT eventid="1422" points="609" swimtime="00:00:26.46" resultid="6797" heatid="10838" lane="6" entrytime="00:00:25.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-13" firstname="Romuald" gender="M" lastname="Kozłowski" nation="POL" athleteid="4343">
              <RESULTS>
                <RESULT eventid="1160" points="331" swimtime="00:00:30.22" resultid="6806" heatid="10695" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1422" points="330" swimtime="00:00:32.44" resultid="6807" heatid="10828" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1638" points="356" swimtime="00:00:37.27" resultid="6808" heatid="10915" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-26" firstname="Tomasz" gender="M" lastname="Wilczęga" nation="POL" athleteid="4349">
              <RESULTS>
                <RESULT eventid="1160" points="456" swimtime="00:00:27.15" resultid="6810" heatid="10689" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-27" firstname="Jan" gender="M" lastname="Peńsko" nation="POL" athleteid="4336">
              <RESULTS>
                <RESULT eventid="1160" points="514" swimtime="00:00:26.10" resultid="6800" heatid="10689" lane="1" />
                <RESULT eventid="1190" points="525" swimtime="00:02:21.26" resultid="6801" heatid="10730" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                    <SPLIT distance="100" swimtime="00:01:04.24" />
                    <SPLIT distance="150" swimtime="00:01:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn w  kat B  30-34  lata" eventid="1332" points="503" swimtime="00:02:20.14" resultid="6802" heatid="10796" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                    <SPLIT distance="100" swimtime="00:01:07.42" />
                    <SPLIT distance="150" swimtime="00:01:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="511" swimtime="00:05:04.83" resultid="6803" heatid="10881" lane="4" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="150" swimtime="00:01:46.96" />
                    <SPLIT distance="200" swimtime="00:02:25.70" />
                    <SPLIT distance="250" swimtime="00:03:10.50" />
                    <SPLIT distance="300" swimtime="00:03:55.61" />
                    <SPLIT distance="350" swimtime="00:04:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="6804" heatid="10892" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="1695" points="451" swimtime="00:04:46.88" resultid="6805" heatid="10935" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:08.67" />
                    <SPLIT distance="150" swimtime="00:01:45.62" />
                    <SPLIT distance="200" swimtime="00:02:23.13" />
                    <SPLIT distance="250" swimtime="00:03:00.43" />
                    <SPLIT distance="300" swimtime="00:03:39.26" />
                    <SPLIT distance="350" swimtime="00:04:16.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="579" swimtime="00:01:52.08" resultid="6818" heatid="10802" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:01:00.09" />
                    <SPLIT distance="150" swimtime="00:01:25.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4336" number="1" />
                    <RELAYPOSITION athleteid="4354" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4330" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4349" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Mężczyzn w  kat B  120-159  lat" eventid="1518" points="671" swimtime="00:01:36.90" resultid="6819" heatid="10872" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.49" />
                    <SPLIT distance="100" swimtime="00:00:48.21" />
                    <SPLIT distance="150" swimtime="00:01:13.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4333" number="1" />
                    <RELAYPOSITION athleteid="4307" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4354" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4330" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1518" status="DNS" swimtime="00:00:00.00" resultid="6820" heatid="10871" lane="5" entrytime="00:01:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MABIA" nation="POL" region="PDL" clubid="4030" name="Masters Białystok">
          <CONTACT email="mbzgloszenia@gmail.com" name="Dominika Michalik" />
          <ATHLETES>
            <ATHLETE birthdate="1966-01-01" firstname="Elżbieta" gender="F" lastname="Piwowarczyk" nation="POL" athleteid="6354">
              <RESULTS>
                <RESULT eventid="1144" points="311" swimtime="00:00:34.99" resultid="6355" heatid="10685" lane="7" entrytime="00:00:34.20" />
                <RESULT eventid="1175" points="271" swimtime="00:03:14.83" resultid="6356" heatid="10715" lane="8" entrytime="00:03:17.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:01:31.86" />
                    <SPLIT distance="150" swimtime="00:02:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="246" swimtime="00:00:43.18" resultid="6357" heatid="10737" lane="9" entrytime="00:00:42.20" />
                <RESULT eventid="1287" points="293" swimtime="00:01:18.38" resultid="6358" heatid="10768" lane="4" entrytime="00:01:17.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="244" swimtime="00:01:32.93" resultid="6359" heatid="10840" lane="5" entrytime="00:01:31.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="270" swimtime="00:02:54.78" resultid="6360" heatid="10853" lane="4" entrytime="00:02:52.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:23.03" />
                    <SPLIT distance="150" swimtime="00:02:09.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="259" swimtime="00:03:14.51" resultid="6361" heatid="10896" lane="9" entrytime="00:03:18.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                    <SPLIT distance="100" swimtime="00:01:35.12" />
                    <SPLIT distance="150" swimtime="00:02:25.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="4031">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat C 35-39 lat" eventid="1113" points="432" swimtime="00:20:24.14" resultid="6337" heatid="10674" lane="4" entrytime="00:20:26.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:01:55.53" />
                    <SPLIT distance="200" swimtime="00:02:36.47" />
                    <SPLIT distance="250" swimtime="00:03:17.25" />
                    <SPLIT distance="300" swimtime="00:03:58.56" />
                    <SPLIT distance="350" swimtime="00:04:39.58" />
                    <SPLIT distance="400" swimtime="00:05:20.72" />
                    <SPLIT distance="450" swimtime="00:06:01.93" />
                    <SPLIT distance="500" swimtime="00:06:43.35" />
                    <SPLIT distance="550" swimtime="00:07:24.60" />
                    <SPLIT distance="600" swimtime="00:08:05.99" />
                    <SPLIT distance="650" swimtime="00:08:46.95" />
                    <SPLIT distance="700" swimtime="00:09:28.06" />
                    <SPLIT distance="750" swimtime="00:10:09.24" />
                    <SPLIT distance="800" swimtime="00:10:50.52" />
                    <SPLIT distance="850" swimtime="00:11:32.41" />
                    <SPLIT distance="900" swimtime="00:12:13.90" />
                    <SPLIT distance="950" swimtime="00:12:55.06" />
                    <SPLIT distance="1000" swimtime="00:13:36.34" />
                    <SPLIT distance="1050" swimtime="00:14:17.15" />
                    <SPLIT distance="1100" swimtime="00:14:57.92" />
                    <SPLIT distance="1150" swimtime="00:15:39.14" />
                    <SPLIT distance="1200" swimtime="00:16:20.44" />
                    <SPLIT distance="1250" swimtime="00:17:02.02" />
                    <SPLIT distance="1300" swimtime="00:17:43.56" />
                    <SPLIT distance="1350" swimtime="00:18:24.86" />
                    <SPLIT distance="1400" swimtime="00:19:05.80" />
                    <SPLIT distance="1450" swimtime="00:19:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="494" swimtime="00:01:05.82" resultid="6338" heatid="10771" lane="0" entrytime="00:01:05.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="347" swimtime="00:00:34.74" resultid="6339" heatid="10823" lane="0" entrytime="00:00:36.15" />
                <RESULT eventid="1467" points="479" swimtime="00:02:24.36" resultid="6340" heatid="10855" lane="7" entrytime="00:02:22.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                    <SPLIT distance="150" swimtime="00:01:46.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="466" swimtime="00:05:04.89" resultid="6341" heatid="10934" lane="6" entrytime="00:05:01.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="150" swimtime="00:01:51.17" />
                    <SPLIT distance="200" swimtime="00:02:30.44" />
                    <SPLIT distance="250" swimtime="00:03:09.64" />
                    <SPLIT distance="300" swimtime="00:03:49.24" />
                    <SPLIT distance="350" swimtime="00:04:28.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Andrzej" gender="M" lastname="Twarowski" nation="POL" athleteid="4037">
              <RESULTS>
                <RESULT eventid="1190" points="179" swimtime="00:03:22.01" resultid="6342" heatid="10722" lane="9" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.88" />
                    <SPLIT distance="100" swimtime="00:01:34.93" />
                    <SPLIT distance="150" swimtime="00:02:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="222" swimtime="00:03:29.61" resultid="6343" heatid="10759" lane="1" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="100" swimtime="00:01:39.65" />
                    <SPLIT distance="150" swimtime="00:02:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="122" swimtime="00:03:44.63" resultid="6344" heatid="10793" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.41" />
                    <SPLIT distance="100" swimtime="00:01:47.54" />
                    <SPLIT distance="150" swimtime="00:02:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="175" swimtime="00:07:15.40" resultid="6345" heatid="10877" lane="3" entrytime="00:07:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.90" />
                    <SPLIT distance="100" swimtime="00:01:46.40" />
                    <SPLIT distance="150" swimtime="00:02:40.54" />
                    <SPLIT distance="200" swimtime="00:03:35.79" />
                    <SPLIT distance="250" swimtime="00:04:35.32" />
                    <SPLIT distance="300" swimtime="00:05:34.40" />
                    <SPLIT distance="350" swimtime="00:06:28.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="182" swimtime="00:03:17.39" resultid="6346" heatid="10901" lane="6" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                    <SPLIT distance="100" swimtime="00:01:33.39" />
                    <SPLIT distance="150" swimtime="00:02:26.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="6347" heatid="10937" lane="4" entrytime="00:06:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Jarosław" gender="M" lastname="Pawlik" nation="POL" athleteid="6348">
              <RESULTS>
                <RESULT eventid="1160" points="192" swimtime="00:00:36.23" resultid="6349" heatid="10695" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="137" swimtime="00:01:30.84" resultid="6350" heatid="10775" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="101" swimtime="00:00:48.15" resultid="6351" heatid="10828" lane="9" entrytime="00:00:42.00" />
                <RESULT eventid="1578" points="62" swimtime="00:02:05.85" resultid="6352" heatid="10886" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="157" swimtime="00:00:48.92" resultid="6353" heatid="10914" lane="4" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="IKMIE" nation="POL" region="PDK" clubid="2877" name="Masters Ikar Mielec">
          <CONTACT city="CHORZELÓW" email="sebastianboicetta@gmail.com" name="SEBASTIAN BOICETTA" phone="501072284" state="PODKA" street="MALINIE 629" zip="39-331" />
          <ATHLETES>
            <ATHLETE birthdate="1988-06-09" firstname="Daniel" gender="M" lastname="Paduch" nation="POL" license="503208700002" athleteid="2878">
              <RESULTS>
                <RESULT eventid="1128" points="464" swimtime="00:18:44.29" resultid="7061" heatid="10679" lane="5" entrytime="00:18:21.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:07.58" />
                    <SPLIT distance="150" swimtime="00:01:43.65" />
                    <SPLIT distance="200" swimtime="00:02:20.10" />
                    <SPLIT distance="250" swimtime="00:02:56.53" />
                    <SPLIT distance="300" swimtime="00:03:33.93" />
                    <SPLIT distance="350" swimtime="00:04:11.19" />
                    <SPLIT distance="400" swimtime="00:04:48.76" />
                    <SPLIT distance="450" swimtime="00:05:26.44" />
                    <SPLIT distance="500" swimtime="00:06:04.47" />
                    <SPLIT distance="550" swimtime="00:06:41.83" />
                    <SPLIT distance="600" swimtime="00:07:20.00" />
                    <SPLIT distance="650" swimtime="00:07:57.63" />
                    <SPLIT distance="700" swimtime="00:08:35.53" />
                    <SPLIT distance="750" swimtime="00:09:13.17" />
                    <SPLIT distance="800" swimtime="00:09:51.57" />
                    <SPLIT distance="850" swimtime="00:10:29.91" />
                    <SPLIT distance="900" swimtime="00:11:07.70" />
                    <SPLIT distance="950" swimtime="00:11:46.47" />
                    <SPLIT distance="1000" swimtime="00:12:24.79" />
                    <SPLIT distance="1050" swimtime="00:13:02.93" />
                    <SPLIT distance="1100" swimtime="00:13:40.99" />
                    <SPLIT distance="1150" swimtime="00:14:19.22" />
                    <SPLIT distance="1200" swimtime="00:14:58.45" />
                    <SPLIT distance="1250" swimtime="00:15:36.45" />
                    <SPLIT distance="1300" swimtime="00:16:14.76" />
                    <SPLIT distance="1350" swimtime="00:16:52.48" />
                    <SPLIT distance="1400" swimtime="00:17:30.53" />
                    <SPLIT distance="1450" swimtime="00:18:07.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="395" swimtime="00:02:35.25" resultid="7062" heatid="10729" lane="2" entrytime="00:02:29.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:02:01.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="505" swimtime="00:02:19.95" resultid="7063" heatid="10796" lane="4" entrytime="00:02:16.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:07.98" />
                    <SPLIT distance="150" swimtime="00:01:44.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="439" swimtime="00:02:14.16" resultid="7064" heatid="10865" lane="7" entrytime="00:02:12.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:07.25" />
                    <SPLIT distance="150" swimtime="00:01:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="401" swimtime="00:05:30.53" resultid="7065" heatid="10881" lane="0" entrytime="00:05:19.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:08.82" />
                    <SPLIT distance="150" swimtime="00:01:57.99" />
                    <SPLIT distance="200" swimtime="00:02:43.88" />
                    <SPLIT distance="250" swimtime="00:03:30.71" />
                    <SPLIT distance="300" swimtime="00:04:18.25" />
                    <SPLIT distance="350" swimtime="00:04:55.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="455" swimtime="00:01:04.75" resultid="7066" heatid="10891" lane="6" entrytime="00:01:03.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="473" swimtime="00:04:42.35" resultid="7067" heatid="10945" lane="2" entrytime="00:04:37.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:08.14" />
                    <SPLIT distance="150" swimtime="00:01:44.12" />
                    <SPLIT distance="200" swimtime="00:02:20.50" />
                    <SPLIT distance="250" swimtime="00:02:56.36" />
                    <SPLIT distance="300" swimtime="00:03:32.33" />
                    <SPLIT distance="350" swimtime="00:04:07.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-24" firstname="Bartek" gender="M" lastname="Kowalik" nation="POL" license="503208700001" athleteid="2886">
              <RESULTS>
                <RESULT eventid="1098" points="319" swimtime="00:11:01.40" resultid="7068" heatid="10673" lane="6" entrytime="00:09:39.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="150" swimtime="00:01:49.05" />
                    <SPLIT distance="200" swimtime="00:02:29.32" />
                    <SPLIT distance="250" swimtime="00:03:10.48" />
                    <SPLIT distance="300" swimtime="00:03:52.20" />
                    <SPLIT distance="350" swimtime="00:04:34.74" />
                    <SPLIT distance="400" swimtime="00:05:17.60" />
                    <SPLIT distance="450" swimtime="00:06:00.49" />
                    <SPLIT distance="500" swimtime="00:06:43.86" />
                    <SPLIT distance="550" swimtime="00:07:27.09" />
                    <SPLIT distance="600" swimtime="00:08:10.89" />
                    <SPLIT distance="650" swimtime="00:08:44.80" />
                    <SPLIT distance="700" swimtime="00:09:37.96" />
                    <SPLIT distance="750" swimtime="00:10:20.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="445" swimtime="00:02:29.27" resultid="7069" heatid="10729" lane="5" entrytime="00:02:26.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="100" swimtime="00:01:10.54" />
                    <SPLIT distance="150" swimtime="00:01:53.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="541" swimtime="00:02:35.83" resultid="7070" heatid="10764" lane="6" entrytime="00:02:36.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:15.73" />
                    <SPLIT distance="150" swimtime="00:01:55.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="522" swimtime="00:01:10.95" resultid="7071" heatid="10819" lane="1" entrytime="00:01:11.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="348" swimtime="00:05:46.63" resultid="7072" heatid="10881" lane="8" entrytime="00:05:14.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:12.41" />
                    <SPLIT distance="150" swimtime="00:02:00.75" />
                    <SPLIT distance="200" swimtime="00:02:46.82" />
                    <SPLIT distance="250" swimtime="00:03:32.68" />
                    <SPLIT distance="300" swimtime="00:04:19.76" />
                    <SPLIT distance="350" swimtime="00:05:04.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="330" swimtime="00:02:41.81" resultid="7073" heatid="10904" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:02:00.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="536" swimtime="00:00:32.51" resultid="7074" heatid="10926" lane="0" entrytime="00:00:31.76" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="7075" heatid="10945" lane="1" entrytime="00:04:39.99" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKRA" nation="POL" region="LBL" clubid="4294" name="Masters Krasnik">
          <CONTACT city="Kraśnik" email="masterskrasnik@gmail.com" internet="www.masterskrasnik.za.pl" name="MIchalczyk Jerzy" phone="601698977" state="LUB" street="Żwirki i Wigury 2" zip="23-204" />
          <ATHLETES>
            <ATHLETE birthdate="1972-11-03" firstname="Agnieszka" gender="F" lastname="Kurzyna" nation="POL" athleteid="4295">
              <RESULTS>
                <RESULT eventid="1226" status="DNS" swimtime="00:00:00.00" resultid="6747" heatid="10735" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1287" status="DNS" swimtime="00:00:00.00" resultid="6748" heatid="10766" lane="7" entrytime="00:01:40.00" />
                <RESULT eventid="1407" status="DNS" swimtime="00:00:00.00" resultid="6749" heatid="10820" lane="4" entrytime="00:00:55.00" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="6750" heatid="10839" lane="3" entrytime="00:02:05.00" />
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="6751" heatid="10894" lane="9" entrytime="00:04:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="4301">
              <RESULTS>
                <RESULT eventid="1242" points="79" swimtime="00:00:55.99" resultid="6752" heatid="10742" lane="7" entrytime="00:00:52.25" />
                <RESULT eventid="1302" points="105" swimtime="00:01:39.27" resultid="6753" heatid="10773" lane="5" entrytime="00:01:42.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="87" swimtime="00:00:50.48" resultid="6754" heatid="10826" lane="5" entrytime="00:00:49.18" />
                <RESULT eventid="1578" points="56" swimtime="00:02:10.05" resultid="6755" heatid="10886" lane="0" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MALUB" nation="POL" region="05" clubid="5645" name="Masters Lublin">
          <CONTACT name="s" />
          <ATHLETES>
            <ATHLETE birthdate="1975-01-01" firstname="Anna" gender="F" lastname="Michalska" nation="POL" athleteid="5655">
              <RESULTS>
                <RESULT eventid="1437" points="359" swimtime="00:01:21.74" resultid="7159" heatid="10842" lane="9" entrytime="00:01:19.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="313" swimtime="00:03:02.57" resultid="7160" heatid="10896" lane="4" entrytime="00:02:57.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:27.31" />
                    <SPLIT distance="150" swimtime="00:02:15.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Konrad" gender="M" lastname="Ćwikła" nation="POL" athleteid="5651">
              <RESULTS>
                <RESULT eventid="1190" points="322" swimtime="00:02:46.24" resultid="7156" heatid="10724" lane="0" entrytime="00:02:55.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:12.82" />
                    <SPLIT distance="150" swimtime="00:02:02.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="430" swimtime="00:01:02.11" resultid="7157" heatid="10781" lane="4" entrytime="00:01:04.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="285" swimtime="00:05:34.28" resultid="7158" heatid="10940" lane="0" entrytime="00:05:59.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:01:17.36" />
                    <SPLIT distance="150" swimtime="00:02:01.09" />
                    <SPLIT distance="200" swimtime="00:02:45.11" />
                    <SPLIT distance="250" swimtime="00:03:29.07" />
                    <SPLIT distance="300" swimtime="00:04:13.06" />
                    <SPLIT distance="350" swimtime="00:04:55.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Rafał" gender="M" lastname="Zielonka" nation="POL" athleteid="5646">
              <RESULTS>
                <RESULT eventid="1098" points="380" swimtime="00:10:23.71" resultid="7152" heatid="10672" lane="4" entrytime="00:10:30.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="150" swimtime="00:01:46.98" />
                    <SPLIT distance="200" swimtime="00:02:25.67" />
                    <SPLIT distance="250" swimtime="00:03:04.29" />
                    <SPLIT distance="300" swimtime="00:03:44.15" />
                    <SPLIT distance="350" swimtime="00:04:23.34" />
                    <SPLIT distance="400" swimtime="00:05:03.03" />
                    <SPLIT distance="450" swimtime="00:05:42.70" />
                    <SPLIT distance="500" swimtime="00:06:22.63" />
                    <SPLIT distance="550" swimtime="00:07:03.14" />
                    <SPLIT distance="600" swimtime="00:07:43.90" />
                    <SPLIT distance="650" swimtime="00:08:24.37" />
                    <SPLIT distance="700" swimtime="00:09:04.90" />
                    <SPLIT distance="750" swimtime="00:09:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="489" swimtime="00:00:59.53" resultid="7153" heatid="10786" lane="6" entrytime="00:00:58.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="489" swimtime="00:02:09.46" resultid="7154" heatid="10865" lane="1" entrytime="00:02:12.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="100" swimtime="00:01:03.80" />
                    <SPLIT distance="150" swimtime="00:01:37.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="482" swimtime="00:04:40.64" resultid="7155" heatid="10944" lane="2" entrytime="00:04:50.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:06.30" />
                    <SPLIT distance="150" swimtime="00:01:41.99" />
                    <SPLIT distance="200" swimtime="00:02:18.21" />
                    <SPLIT distance="250" swimtime="00:02:54.25" />
                    <SPLIT distance="300" swimtime="00:03:30.28" />
                    <SPLIT distance="350" swimtime="00:04:06.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MABIAL" nation="POL" region="PDL" clubid="4007" name="Masters Team Biała Podlaska">
          <CONTACT internet="wilhelmg@poczta.onet.pl" name="Gromisz" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-15" firstname="Michał" gender="M" lastname="Jagiełło" nation="POL" athleteid="4026">
              <RESULTS>
                <RESULT eventid="1160" points="635" swimtime="00:00:24.32" resultid="6330" heatid="10711" lane="8" entrytime="00:00:24.64" />
                <RESULT eventid="1302" points="597" swimtime="00:00:55.71" resultid="6331" heatid="10787" lane="6" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="522" swimtime="00:00:27.84" resultid="6332" heatid="10837" lane="2" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-07" firstname="Robert" gender="M" lastname="Jagiełło" nation="POL" athleteid="4023">
              <RESULTS>
                <RESULT eventid="1160" points="194" swimtime="00:00:36.11" resultid="6328" heatid="10696" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1392" points="154" swimtime="00:01:46.50" resultid="6329" heatid="10812" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-12-27" firstname="Renata" gender="F" lastname="Kasprowicz" nation="POL" athleteid="4008">
              <RESULTS>
                <RESULT eventid="1144" points="454" swimtime="00:00:30.87" resultid="6315" heatid="10687" lane="2" entrytime="00:00:30.35" />
                <RESULT eventid="1257" points="355" swimtime="00:03:16.41" resultid="6316" heatid="10756" lane="9" entrytime="00:03:09.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.61" />
                    <SPLIT distance="100" swimtime="00:01:33.68" />
                    <SPLIT distance="150" swimtime="00:02:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="392" swimtime="00:01:27.87" resultid="6317" heatid="10808" lane="7" entrytime="00:01:24.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="369" swimtime="00:00:34.05" resultid="6318" heatid="10823" lane="4" entrytime="00:00:33.54" />
                <RESULT eventid="1623" points="417" swimtime="00:00:39.44" resultid="6319" heatid="10911" lane="0" entrytime="00:00:38.51" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Iga" gender="F" lastname="Olszanowska" nation="POL" athleteid="4014">
              <RESULTS>
                <RESULT eventid="1144" points="471" swimtime="00:00:30.49" resultid="6320" heatid="10688" lane="8" entrytime="00:00:29.30" />
                <RESULT eventid="1175" points="389" swimtime="00:02:52.72" resultid="6321" heatid="10718" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:20.46" />
                    <SPLIT distance="150" swimtime="00:02:10.42" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat C  35-39  lat" eventid="1226" points="480" swimtime="00:00:34.56" resultid="6322" heatid="10739" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1287" points="468" swimtime="00:01:07.05" resultid="6323" heatid="10771" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="389" swimtime="00:01:28.15" resultid="6324" heatid="10808" lane="3" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="341" swimtime="00:06:21.07" resultid="6325" heatid="10875" lane="1" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:02:14.34" />
                    <SPLIT distance="200" swimtime="00:03:05.30" />
                    <SPLIT distance="250" swimtime="00:03:57.74" />
                    <SPLIT distance="300" swimtime="00:04:52.18" />
                    <SPLIT distance="350" swimtime="00:05:38.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="374" swimtime="00:01:16.98" resultid="6326" heatid="10884" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="392" swimtime="00:00:40.27" resultid="6327" heatid="10911" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WIKRA" nation="POL" region="MAL" clubid="3180" name="Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Tomasz Doniec" phone="693703490" />
          <ATHLETES>
            <ATHLETE birthdate="1978-09-30" firstname="Szymon" gender="M" lastname="Łenyk" nation="POL" athleteid="3270">
              <RESULTS>
                <RESULT eventid="1160" points="171" swimtime="00:00:37.64" resultid="3271" heatid="10694" lane="8" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1190" points="96" swimtime="00:04:08.66" resultid="3272" heatid="10719" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.97" />
                    <SPLIT distance="100" swimtime="00:02:01.92" />
                    <SPLIT distance="150" swimtime="00:03:07.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="103" swimtime="00:00:51.21" resultid="3273" heatid="10743" lane="8" entrytime="00:00:50.00" entrycourse="LCM" />
                <RESULT eventid="1302" points="141" swimtime="00:01:30.11" resultid="3274" heatid="10775" lane="7" entrytime="00:01:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="141" swimtime="00:01:49.59" resultid="3275" heatid="10811" lane="9" entrytime="00:01:48.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="3276" heatid="10856" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Karolina" gender="F" lastname="Górka" nation="POL" athleteid="3306">
              <RESULTS>
                <RESULT eventid="1144" points="401" swimtime="00:00:32.17" resultid="3307" heatid="10687" lane="9" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1257" points="342" swimtime="00:03:18.87" resultid="3308" heatid="10755" lane="1" entrytime="00:03:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                    <SPLIT distance="100" swimtime="00:01:34.35" />
                    <SPLIT distance="150" swimtime="00:02:26.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="342" swimtime="00:01:14.39" resultid="3309" heatid="10769" lane="2" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="356" swimtime="00:01:30.73" resultid="3310" heatid="10807" lane="9" entrytime="00:01:35.00" entrycourse="LCM" />
                <RESULT eventid="1467" points="272" swimtime="00:02:54.26" resultid="3311" heatid="10854" lane="9" entrytime="00:02:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                    <SPLIT distance="100" swimtime="00:01:23.34" />
                    <SPLIT distance="150" swimtime="00:02:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="396" swimtime="00:00:40.12" resultid="3312" heatid="10909" lane="3" entrytime="00:00:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-26" firstname="Iwona" gender="F" lastname="Bednarczyk" nation="POL" athleteid="3200">
              <RESULTS>
                <RESULT eventid="1059" points="88" swimtime="00:18:09.65" resultid="3201" heatid="10666" lane="8" entrytime="00:18:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.73" />
                    <SPLIT distance="100" swimtime="00:01:59.68" />
                    <SPLIT distance="150" swimtime="00:03:08.32" />
                    <SPLIT distance="200" swimtime="00:04:16.31" />
                    <SPLIT distance="250" swimtime="00:05:25.56" />
                    <SPLIT distance="300" swimtime="00:06:34.42" />
                    <SPLIT distance="350" swimtime="00:07:43.73" />
                    <SPLIT distance="400" swimtime="00:08:55.45" />
                    <SPLIT distance="450" swimtime="00:10:03.31" />
                    <SPLIT distance="500" swimtime="00:11:12.65" />
                    <SPLIT distance="550" swimtime="00:12:21.43" />
                    <SPLIT distance="600" swimtime="00:13:31.23" />
                    <SPLIT distance="650" swimtime="00:14:41.02" />
                    <SPLIT distance="700" swimtime="00:15:51.46" />
                    <SPLIT distance="750" swimtime="00:17:02.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="85" swimtime="00:04:46.01" resultid="3202" heatid="10713" lane="9" entrytime="00:04:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.11" />
                    <SPLIT distance="100" swimtime="00:02:23.42" />
                    <SPLIT distance="150" swimtime="00:03:43.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="68" swimtime="00:01:06.00" resultid="3203" heatid="10735" lane="0" entrytime="00:00:59.00" entrycourse="LCM" />
                <RESULT eventid="1287" points="94" swimtime="00:01:54.37" resultid="3204" heatid="10766" lane="0" entrytime="00:01:50.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="57" swimtime="00:01:03.23" resultid="3205" heatid="10820" lane="2" entrytime="00:01:02.00" entrycourse="LCM" />
                <RESULT eventid="1467" points="98" swimtime="00:04:04.70" resultid="3206" heatid="10851" lane="6" entrytime="00:04:13.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.70" />
                    <SPLIT distance="100" swimtime="00:01:55.52" />
                    <SPLIT distance="150" swimtime="00:03:00.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="57" swimtime="00:02:23.90" resultid="3207" heatid="10882" lane="4" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="86" swimtime="00:08:53.65" resultid="3208" heatid="10931" lane="8" entrytime="00:08:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.11" />
                    <SPLIT distance="100" swimtime="00:01:55.82" />
                    <SPLIT distance="150" swimtime="00:03:04.58" />
                    <SPLIT distance="200" swimtime="00:04:16.07" />
                    <SPLIT distance="250" swimtime="00:05:26.97" />
                    <SPLIT distance="300" swimtime="00:06:37.59" />
                    <SPLIT distance="350" swimtime="00:07:45.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-11-06" firstname="Małgorzata" gender="F" lastname="Wach" nation="POL" athleteid="3256">
              <RESULTS>
                <RESULT eventid="1144" points="232" swimtime="00:00:38.61" resultid="3257" heatid="10684" lane="9" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1226" points="264" swimtime="00:00:42.14" resultid="3258" heatid="10737" lane="8" entrytime="00:00:42.00" entrycourse="LCM" />
                <RESULT eventid="1287" points="238" swimtime="00:01:23.94" resultid="3259" heatid="10767" lane="5" entrytime="00:01:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="220" swimtime="00:01:36.24" resultid="3260" heatid="10840" lane="4" entrytime="00:01:31.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="208" swimtime="00:03:10.63" resultid="3261" heatid="10853" lane="0" entrytime="00:03:07.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                    <SPLIT distance="100" swimtime="00:01:31.16" />
                    <SPLIT distance="150" swimtime="00:02:21.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="3262" heatid="10895" lane="2" entrytime="00:03:25.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-04" firstname="Małgorzata" gender="F" lastname="Skalska" nation="POL" athleteid="3283">
              <RESULTS>
                <RESULT eventid="1175" points="163" swimtime="00:03:50.76" resultid="3284" heatid="10712" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.92" />
                    <SPLIT distance="100" swimtime="00:01:56.60" />
                    <SPLIT distance="150" swimtime="00:02:56.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="199" swimtime="00:03:58.09" resultid="3285" heatid="10755" lane="9" entrytime="00:03:34.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.79" />
                    <SPLIT distance="100" swimtime="00:01:51.11" />
                    <SPLIT distance="150" swimtime="00:02:55.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="192" swimtime="00:01:30.20" resultid="3286" heatid="10767" lane="2" entrytime="00:01:27.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="197" swimtime="00:01:50.51" resultid="3287" heatid="10805" lane="7" entrytime="00:01:44.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="3288" heatid="10852" lane="3" entrytime="00:03:20.50" entrycourse="LCM" />
                <RESULT eventid="1674" points="159" swimtime="00:07:15.88" resultid="3289" heatid="10932" lane="7" entrytime="00:07:07.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.58" />
                    <SPLIT distance="100" swimtime="00:01:42.17" />
                    <SPLIT distance="150" swimtime="00:02:38.39" />
                    <SPLIT distance="200" swimtime="00:03:35.82" />
                    <SPLIT distance="250" swimtime="00:04:32.46" />
                    <SPLIT distance="300" swimtime="00:05:29.19" />
                    <SPLIT distance="350" swimtime="00:06:24.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="3263">
              <RESULTS>
                <RESULT eventid="1226" points="109" swimtime="00:00:56.52" resultid="3264" heatid="10735" lane="7" entrytime="00:00:56.00" entrycourse="LCM" />
                <RESULT eventid="1257" points="142" swimtime="00:04:26.61" resultid="3265" heatid="10753" lane="7" entrytime="00:04:39.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.04" />
                    <SPLIT distance="100" swimtime="00:02:12.50" />
                    <SPLIT distance="150" swimtime="00:03:20.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="123" swimtime="00:02:09.13" resultid="3266" heatid="10804" lane="0" entrytime="00:02:09.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="108" swimtime="00:02:01.93" resultid="3267" heatid="10840" lane="9" entrytime="00:01:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="115" swimtime="00:04:14.44" resultid="3268" heatid="10894" lane="1" entrytime="00:04:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.75" />
                    <SPLIT distance="100" swimtime="00:02:06.45" />
                    <SPLIT distance="150" swimtime="00:03:10.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="115" swimtime="00:01:00.52" resultid="3269" heatid="10905" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-03-06" firstname="Ewa" gender="F" lastname="Rupp" nation="POL" athleteid="3211">
              <RESULTS>
                <RESULT eventid="1144" points="139" swimtime="00:00:45.74" resultid="3212" heatid="10682" lane="0" entrytime="00:00:47.40" entrycourse="LCM" />
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="3213" heatid="10713" lane="0" entrytime="00:04:35.00" entrycourse="LCM" />
                <RESULT eventid="1226" points="116" swimtime="00:00:55.37" resultid="3214" heatid="10735" lane="8" entrytime="00:00:56.50" entrycourse="LCM" />
                <RESULT eventid="1287" points="106" swimtime="00:01:49.97" resultid="3215" heatid="10766" lane="9" entrytime="00:01:53.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" status="DNS" swimtime="00:00:00.00" resultid="3216" heatid="10820" lane="3" entrytime="00:00:59.90" entrycourse="LCM" />
                <RESULT eventid="1437" points="94" swimtime="00:02:07.59" resultid="3217" heatid="10839" lane="6" entrytime="00:02:09.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="62" swimtime="00:02:19.80" resultid="3218" heatid="10882" lane="5" entrytime="00:02:35.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="99" swimtime="00:04:27.76" resultid="3219" heatid="10894" lane="8" entrytime="00:04:35.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.13" />
                    <SPLIT distance="100" swimtime="00:02:12.58" />
                    <SPLIT distance="150" swimtime="00:03:22.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-03-22" firstname="Sandra" gender="F" lastname="Wolska" nation="POL" athleteid="3190">
              <RESULTS>
                <RESULT eventid="1059" points="230" swimtime="00:13:10.36" resultid="3191" heatid="10665" lane="2" />
                <RESULT eventid="1144" points="346" swimtime="00:00:33.80" resultid="3192" heatid="10686" lane="9" entrytime="00:00:33.58" entrycourse="LCM" />
                <RESULT eventid="1175" points="267" swimtime="00:03:15.71" resultid="3193" heatid="10715" lane="3" entrytime="00:03:11.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                    <SPLIT distance="100" swimtime="00:01:38.75" />
                    <SPLIT distance="150" swimtime="00:02:30.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="310" swimtime="00:03:25.34" resultid="3194" heatid="10755" lane="6" entrytime="00:03:19.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.91" />
                    <SPLIT distance="100" swimtime="00:01:36.83" />
                    <SPLIT distance="150" swimtime="00:02:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1317" points="230" swimtime="00:03:18.79" resultid="3195" heatid="10790" lane="8" entrytime="00:03:41.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                    <SPLIT distance="100" swimtime="00:01:31.46" />
                    <SPLIT distance="150" swimtime="00:02:24.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="324" swimtime="00:01:33.64" resultid="3196" heatid="10807" lane="3" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="288" swimtime="00:06:43.08" resultid="3197" heatid="10874" lane="7" entrytime="00:06:53.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:31.65" />
                    <SPLIT distance="150" swimtime="00:02:27.86" />
                    <SPLIT distance="200" swimtime="00:03:23.08" />
                    <SPLIT distance="250" swimtime="00:04:15.91" />
                    <SPLIT distance="300" swimtime="00:05:09.80" />
                    <SPLIT distance="350" swimtime="00:05:57.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="244" swimtime="00:03:18.47" resultid="3198" heatid="10895" lane="1" entrytime="00:03:26.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.28" />
                    <SPLIT distance="100" swimtime="00:01:35.03" />
                    <SPLIT distance="150" swimtime="00:02:26.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="392" swimtime="00:00:40.26" resultid="3199" heatid="10909" lane="4" entrytime="00:00:41.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" athleteid="3220">
              <RESULTS>
                <RESULT eventid="1144" points="574" swimtime="00:00:28.55" resultid="3221" heatid="10688" lane="3" entrytime="00:00:27.60" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat A  25-29 lat" eventid="1175" points="621" swimtime="00:02:27.78" resultid="3222" heatid="10718" lane="4" entrytime="00:02:26.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                    <SPLIT distance="100" swimtime="00:01:11.27" />
                    <SPLIT distance="150" swimtime="00:01:53.82" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat A  25-29  lat" eventid="1257" points="586" swimtime="00:02:46.20" resultid="3223" heatid="10756" lane="5" entrytime="00:02:48.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="100" swimtime="00:01:20.22" />
                    <SPLIT distance="150" swimtime="00:02:03.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="610" swimtime="00:01:01.37" resultid="3224" heatid="10771" lane="3" entrytime="00:01:00.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat A  25-29  lat" eventid="1467" points="642" swimtime="00:02:10.92" resultid="3225" heatid="10855" lane="4" entrytime="00:02:11.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:01:04.19" />
                    <SPLIT distance="150" swimtime="00:01:38.26" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat A  25-29  lat" eventid="1525" points="618" swimtime="00:05:12.56" resultid="3226" heatid="10875" lane="4" entrytime="00:05:14.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:11.51" />
                    <SPLIT distance="150" swimtime="00:01:53.22" />
                    <SPLIT distance="200" swimtime="00:02:33.67" />
                    <SPLIT distance="250" swimtime="00:03:17.54" />
                    <SPLIT distance="300" swimtime="00:04:01.24" />
                    <SPLIT distance="350" swimtime="00:04:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="590" swimtime="00:00:35.13" resultid="3227" heatid="10911" lane="4" entrytime="00:00:35.12" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1674" points="588" swimtime="00:04:42.13" resultid="3228" heatid="10934" lane="4" entrytime="00:04:38.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:01:08.13" />
                    <SPLIT distance="150" swimtime="00:01:45.00" />
                    <SPLIT distance="200" swimtime="00:02:21.72" />
                    <SPLIT distance="250" swimtime="00:02:58.31" />
                    <SPLIT distance="300" swimtime="00:03:34.29" />
                    <SPLIT distance="350" swimtime="00:04:09.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-25" firstname="Agnieszka" gender="F" lastname="Krupa" nation="POL" athleteid="3234">
              <RESULTS>
                <RESULT eventid="1059" status="DNF" swimtime="00:00:00.00" resultid="3235" heatid="10665" lane="6" />
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="3236" heatid="10682" lane="5" entrytime="00:00:42.46" entrycourse="LCM" />
                <RESULT eventid="1226" points="153" swimtime="00:00:50.58" resultid="3237" heatid="10735" lane="6" entrytime="00:00:51.12" entrycourse="LCM" />
                <RESULT eventid="1287" points="164" swimtime="00:01:34.92" resultid="3238" heatid="10767" lane="9" entrytime="00:01:31.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="153" swimtime="00:03:31.04" resultid="3239" heatid="10852" lane="6" entrytime="00:03:26.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                    <SPLIT distance="100" swimtime="00:01:39.77" />
                    <SPLIT distance="150" swimtime="00:02:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" status="DNS" swimtime="00:00:00.00" resultid="3240" heatid="10930" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-25" firstname="Jerzy" gender="M" lastname="Korba" nation="POL" athleteid="3290">
              <RESULTS>
                <RESULT eventid="1098" points="358" swimtime="00:10:36.33" resultid="3291" heatid="10673" lane="0" entrytime="00:10:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:10.97" />
                    <SPLIT distance="150" swimtime="00:01:49.42" />
                    <SPLIT distance="200" swimtime="00:02:28.72" />
                    <SPLIT distance="250" swimtime="00:03:08.54" />
                    <SPLIT distance="300" swimtime="00:03:48.85" />
                    <SPLIT distance="350" swimtime="00:04:29.19" />
                    <SPLIT distance="400" swimtime="00:05:09.71" />
                    <SPLIT distance="450" swimtime="00:05:50.29" />
                    <SPLIT distance="500" swimtime="00:06:31.13" />
                    <SPLIT distance="550" swimtime="00:07:12.27" />
                    <SPLIT distance="600" swimtime="00:07:53.41" />
                    <SPLIT distance="650" swimtime="00:08:35.05" />
                    <SPLIT distance="700" swimtime="00:09:16.44" />
                    <SPLIT distance="750" swimtime="00:09:57.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="413" swimtime="00:00:28.07" resultid="3292" heatid="10706" lane="4" entrytime="00:00:27.46" entrycourse="LCM" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="3293" heatid="10727" lane="5" entrytime="00:02:37.40" entrycourse="LCM" />
                <RESULT eventid="1272" points="345" swimtime="00:03:00.93" resultid="3294" heatid="10757" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:01:27.81" />
                    <SPLIT distance="150" swimtime="00:02:16.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="3295" heatid="10784" lane="4" entrytime="00:01:00.50" entrycourse="LCM" />
                <RESULT eventid="1392" points="376" swimtime="00:01:19.09" resultid="3296" heatid="10817" lane="1" entrytime="00:01:18.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="3297" heatid="10864" lane="7" entrytime="00:02:15.00" entrycourse="LCM" />
                <RESULT eventid="1638" points="437" swimtime="00:00:34.80" resultid="3298" heatid="10924" lane="2" entrytime="00:00:33.96" entrycourse="LCM" />
                <RESULT eventid="1695" points="343" swimtime="00:05:14.21" resultid="3299" heatid="10943" lane="5" entrytime="00:05:00.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:01:54.78" />
                    <SPLIT distance="200" swimtime="00:02:35.14" />
                    <SPLIT distance="250" swimtime="00:03:15.55" />
                    <SPLIT distance="300" swimtime="00:03:55.75" />
                    <SPLIT distance="350" swimtime="00:04:36.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-16" firstname="Tomasz" gender="M" lastname="Doniec" nation="POL" athleteid="3181">
              <RESULTS>
                <RESULT eventid="1272" points="212" swimtime="00:03:32.76" resultid="3182" heatid="10759" lane="3" entrytime="00:03:28.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                    <SPLIT distance="100" swimtime="00:01:45.63" />
                    <SPLIT distance="150" swimtime="00:02:43.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="257" swimtime="00:01:29.75" resultid="3183" heatid="10813" lane="6" entrytime="00:01:30.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="323" swimtime="00:00:38.48" resultid="3184" heatid="10920" lane="8" entrytime="00:00:38.08" entrycourse="LCM" />
                <RESULT eventid="1695" points="132" swimtime="00:07:12.08" resultid="3185" heatid="10937" lane="7" entrytime="00:06:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.35" />
                    <SPLIT distance="100" swimtime="00:01:42.17" />
                    <SPLIT distance="150" swimtime="00:02:39.33" />
                    <SPLIT distance="200" swimtime="00:03:35.75" />
                    <SPLIT distance="250" swimtime="00:04:31.80" />
                    <SPLIT distance="300" swimtime="00:05:29.69" />
                    <SPLIT distance="350" swimtime="00:06:23.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1930-05-04" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="3241">
              <RESULTS>
                <RESULT eventid="1160" points="105" swimtime="00:00:44.27" resultid="3242" heatid="10691" lane="4" entrytime="00:00:44.00" entrycourse="LCM" />
                <RESULT eventid="1190" points="60" swimtime="00:04:50.83" resultid="3243" heatid="10720" lane="8" entrytime="00:04:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.51" />
                    <SPLIT distance="100" swimtime="00:02:34.23" />
                    <SPLIT distance="150" swimtime="00:03:52.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="69" swimtime="00:00:58.40" resultid="3244" heatid="10741" lane="1" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="1302" points="80" swimtime="00:01:48.59" resultid="3245" heatid="10773" lane="4" entrytime="00:01:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="68" swimtime="00:02:19.34" resultid="3246" heatid="10810" lane="0" entrytime="00:02:02.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="70" swimtime="00:04:06.62" resultid="3247" heatid="10857" lane="0" entrytime="00:04:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.94" />
                    <SPLIT distance="100" swimtime="00:01:56.02" />
                    <SPLIT distance="150" swimtime="00:03:00.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="85" swimtime="00:00:59.96" resultid="3248" heatid="10913" lane="7" entrytime="00:01:00.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-22" firstname="Mateusz" gender="M" lastname="Dybek" nation="POL" athleteid="3186">
              <RESULTS>
                <RESULT eventid="1128" points="336" swimtime="00:20:52.53" resultid="3187" heatid="10678" lane="6" entrytime="00:21:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                    <SPLIT distance="100" swimtime="00:01:14.41" />
                    <SPLIT distance="150" swimtime="00:01:55.43" />
                    <SPLIT distance="200" swimtime="00:02:36.77" />
                    <SPLIT distance="250" swimtime="00:03:18.34" />
                    <SPLIT distance="300" swimtime="00:04:00.45" />
                    <SPLIT distance="350" swimtime="00:04:42.23" />
                    <SPLIT distance="400" swimtime="00:05:24.53" />
                    <SPLIT distance="450" swimtime="00:06:06.76" />
                    <SPLIT distance="500" swimtime="00:06:49.52" />
                    <SPLIT distance="550" swimtime="00:07:32.12" />
                    <SPLIT distance="600" swimtime="00:08:14.81" />
                    <SPLIT distance="650" swimtime="00:08:56.77" />
                    <SPLIT distance="700" swimtime="00:09:39.45" />
                    <SPLIT distance="750" swimtime="00:10:21.16" />
                    <SPLIT distance="800" swimtime="00:11:03.35" />
                    <SPLIT distance="850" swimtime="00:11:45.00" />
                    <SPLIT distance="900" swimtime="00:12:27.75" />
                    <SPLIT distance="950" swimtime="00:13:10.25" />
                    <SPLIT distance="1000" swimtime="00:13:52.55" />
                    <SPLIT distance="1050" swimtime="00:14:34.45" />
                    <SPLIT distance="1100" swimtime="00:15:16.83" />
                    <SPLIT distance="1150" swimtime="00:15:58.84" />
                    <SPLIT distance="1200" swimtime="00:16:41.30" />
                    <SPLIT distance="1250" swimtime="00:17:23.54" />
                    <SPLIT distance="1300" swimtime="00:18:06.28" />
                    <SPLIT distance="1350" swimtime="00:18:48.81" />
                    <SPLIT distance="1400" swimtime="00:19:30.97" />
                    <SPLIT distance="1450" swimtime="00:20:12.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="436" swimtime="00:00:27.56" resultid="3188" heatid="10708" lane="7" entrytime="00:00:26.60" entrycourse="LCM" />
                <RESULT eventid="1302" points="467" swimtime="00:01:00.43" resultid="3189" heatid="10786" lane="1" entrytime="00:00:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-12" firstname="Janusz" gender="M" lastname="Mrozik" nation="POL" athleteid="3229">
              <RESULTS>
                <RESULT eventid="1272" points="60" swimtime="00:05:22.76" resultid="3230" heatid="10757" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.69" />
                    <SPLIT distance="100" swimtime="00:02:40.57" />
                    <SPLIT distance="150" swimtime="00:04:03.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="51" swimtime="00:02:33.96" resultid="3231" heatid="10809" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="51" swimtime="00:04:34.05" resultid="3232" heatid="10856" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.09" />
                    <SPLIT distance="100" swimtime="00:02:14.03" />
                    <SPLIT distance="150" swimtime="00:03:25.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="47" swimtime="00:01:13.20" resultid="3233" heatid="10912" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-19" firstname="Paullina" gender="F" lastname="Palka" nation="POL" athleteid="3209">
              <RESULTS>
                <RESULT eventid="1593" points="328" swimtime="00:02:59.89" resultid="3210" heatid="10897" lane="9" entrytime="00:02:55.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                    <SPLIT distance="150" swimtime="00:02:14.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-02-07" firstname="Bogdan" gender="M" lastname="Szczurek" nation="POL" athleteid="3277">
              <RESULTS>
                <RESULT eventid="1242" points="65" swimtime="00:00:59.50" resultid="3278" heatid="10740" lane="3" />
                <RESULT eventid="1302" points="56" swimtime="00:02:02.26" resultid="3279" heatid="10772" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="52" swimtime="00:02:18.81" resultid="3280" heatid="10843" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="54" swimtime="00:04:29.43" resultid="3281" heatid="10856" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.37" />
                    <SPLIT distance="100" swimtime="00:02:05.76" />
                    <SPLIT distance="150" swimtime="00:03:17.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="52" swimtime="00:04:59.45" resultid="3282" heatid="10898" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.98" />
                    <SPLIT distance="100" swimtime="00:02:27.89" />
                    <SPLIT distance="150" swimtime="00:03:47.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-10" firstname="Dariusz" gender="M" lastname="Wesołowski" nation="POL" athleteid="3300">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="3301" heatid="10704" lane="5" entrytime="00:00:28.20" entrycourse="LCM" />
                <RESULT eventid="1242" points="166" swimtime="00:00:43.71" resultid="3302" heatid="10743" lane="9" entrytime="00:00:50.00" entrycourse="LCM" />
                <RESULT eventid="1302" points="311" swimtime="00:01:09.18" resultid="3303" heatid="10781" lane="0" entrytime="00:01:06.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="318" swimtime="00:00:32.83" resultid="3304" heatid="10831" lane="7" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1482" points="228" swimtime="00:02:46.90" resultid="3305" heatid="10860" lane="5" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:18.69" />
                    <SPLIT distance="150" swimtime="00:02:04.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-01" firstname="Grzegorz" gender="M" lastname="Grzybczyk" nation="POL" athleteid="3249">
              <RESULTS>
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="3250" heatid="10742" lane="2" entrytime="00:00:52.00" entrycourse="LCM" />
                <RESULT eventid="1272" points="92" swimtime="00:04:41.28" resultid="3251" heatid="10758" lane="9" entrytime="00:04:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.57" />
                    <SPLIT distance="100" swimtime="00:02:12.70" />
                    <SPLIT distance="150" swimtime="00:03:26.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="85" swimtime="00:02:09.81" resultid="3252" heatid="10810" lane="1" entrytime="00:02:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="58" swimtime="00:02:13.68" resultid="3253" heatid="10844" lane="3" entrytime="00:02:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="47" swimtime="00:02:17.40" resultid="3254" heatid="10885" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="91" swimtime="00:00:58.58" resultid="3255" heatid="10913" lane="3" entrytime="00:00:56.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" name="Wisła 4" number="4">
              <RESULTS>
                <RESULT eventid="1368" points="200" swimtime="00:02:39.57" resultid="3315" heatid="10800" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.41" />
                    <SPLIT distance="150" swimtime="00:01:24.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3249" number="1" />
                    <RELAYPOSITION athleteid="3181" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3300" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3290" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" name="Wisła 5" number="5">
              <RESULTS>
                <RESULT eventid="1368" points="63" swimtime="00:03:54.15" resultid="3316" heatid="10799" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.33" />
                    <SPLIT distance="100" swimtime="00:02:14.93" />
                    <SPLIT distance="150" swimtime="00:03:06.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3277" number="1" />
                    <RELAYPOSITION athleteid="3229" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3270" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3241" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F" name="Wisła 3" number="3">
              <RESULTS>
                <RESULT eventid="1347" points="142" swimtime="00:03:23.38" resultid="3314" heatid="10797" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.13" />
                    <SPLIT distance="100" swimtime="00:01:44.20" />
                    <SPLIT distance="150" swimtime="00:02:47.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3263" number="1" />
                    <RELAYPOSITION athleteid="3283" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3211" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3256" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" name="Wisła 1" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:49.41" resultid="3313" heatid="10731" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                    <SPLIT distance="100" swimtime="00:01:21.07" />
                    <SPLIT distance="150" swimtime="00:02:11.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3211" number="1" />
                    <RELAYPOSITION athleteid="3181" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3200" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3270" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="Wisła 6" number="6">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:52.62" resultid="3317" heatid="10927" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="150" swimtime="00:02:13.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3209" number="1" />
                    <RELAYPOSITION athleteid="3181" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3249" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3283" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" name="Wisła 7" number="7">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:03:40.60" resultid="3318" heatid="10927" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.78" />
                    <SPLIT distance="100" swimtime="00:02:02.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3277" number="1" />
                    <RELAYPOSITION athleteid="3263" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3234" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3241" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAZDZ" nation="POL" region="OPO" clubid="6074" name="MASTERS Zdzieszowice">
          <CONTACT email="masters.zdzieszowice@gmail.com" name="Jajuga" phone="505127695" />
          <ATHLETES>
            <ATHLETE birthdate="1980-01-26" firstname="Katarzyna" gender="F" lastname="Gniot" nation="POL" athleteid="6099">
              <RESULTS>
                <RESULT eventid="1144" points="240" swimtime="00:00:38.17" resultid="8848" heatid="10684" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1175" points="150" swimtime="00:03:57.11" resultid="8849" heatid="10713" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.18" />
                    <SPLIT distance="100" swimtime="00:02:00.90" />
                    <SPLIT distance="150" swimtime="00:03:05.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="136" swimtime="00:00:52.60" resultid="8850" heatid="10735" lane="2" entrytime="00:00:55.00" />
                <RESULT eventid="1257" points="177" swimtime="00:04:07.64" resultid="8851" heatid="10754" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.00" />
                    <SPLIT distance="100" swimtime="00:02:01.19" />
                    <SPLIT distance="150" swimtime="00:03:05.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="169" swimtime="00:01:56.23" resultid="8852" heatid="10804" lane="6" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="124" swimtime="00:01:56.37" resultid="8853" heatid="10839" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="129" swimtime="00:04:04.98" resultid="8854" heatid="10894" lane="2" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.12" />
                    <SPLIT distance="100" swimtime="00:02:02.03" />
                    <SPLIT distance="150" swimtime="00:03:04.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="184" swimtime="00:00:51.83" resultid="8855" heatid="10907" lane="0" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-23" firstname="Ewelina" gender="F" lastname="Cuch" nation="POL" athleteid="6108" />
            <ATHLETE birthdate="1986-02-15" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="6081">
              <RESULTS>
                <RESULT eventid="1098" points="404" swimtime="00:10:11.44" resultid="8832" heatid="10672" lane="1" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                    <SPLIT distance="150" swimtime="00:01:50.20" />
                    <SPLIT distance="200" swimtime="00:02:29.29" />
                    <SPLIT distance="250" swimtime="00:03:07.86" />
                    <SPLIT distance="300" swimtime="00:03:46.71" />
                    <SPLIT distance="350" swimtime="00:04:25.11" />
                    <SPLIT distance="400" swimtime="00:05:03.78" />
                    <SPLIT distance="450" swimtime="00:05:42.33" />
                    <SPLIT distance="500" swimtime="00:06:21.59" />
                    <SPLIT distance="550" swimtime="00:07:00.77" />
                    <SPLIT distance="600" swimtime="00:07:39.75" />
                    <SPLIT distance="650" swimtime="00:08:17.74" />
                    <SPLIT distance="700" swimtime="00:08:56.18" />
                    <SPLIT distance="750" swimtime="00:09:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="487" swimtime="00:02:24.82" resultid="8833" heatid="10730" lane="0" entrytime="00:02:25.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                    <SPLIT distance="100" swimtime="00:01:07.22" />
                    <SPLIT distance="150" swimtime="00:01:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="8834" heatid="10785" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="1332" points="428" swimtime="00:02:27.91" resultid="8835" heatid="10796" lane="2" entrytime="00:02:26.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="464" swimtime="00:02:11.74" resultid="8836" heatid="10865" lane="2" entrytime="00:02:12.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                    <SPLIT distance="100" swimtime="00:01:04.22" />
                    <SPLIT distance="150" swimtime="00:01:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="468" swimtime="00:05:13.87" resultid="8837" heatid="10881" lane="7" entrytime="00:05:12.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:01:11.35" />
                    <SPLIT distance="150" swimtime="00:01:54.09" />
                    <SPLIT distance="200" swimtime="00:02:35.96" />
                    <SPLIT distance="250" swimtime="00:03:20.45" />
                    <SPLIT distance="300" swimtime="00:04:04.28" />
                    <SPLIT distance="350" swimtime="00:04:39.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="513" swimtime="00:01:02.21" resultid="8838" heatid="10891" lane="3" entrytime="00:01:01.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="8839" heatid="10945" lane="9" entrytime="00:04:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-18" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="6075">
              <RESULTS>
                <RESULT eventid="1175" points="328" swimtime="00:03:02.74" resultid="8827" heatid="10716" lane="3" entrytime="00:03:01.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:26.37" />
                    <SPLIT distance="150" swimtime="00:02:20.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1317" points="245" swimtime="00:03:14.57" resultid="8828" heatid="10790" lane="3" entrytime="00:03:11.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.87" />
                    <SPLIT distance="100" swimtime="00:01:35.19" />
                    <SPLIT distance="150" swimtime="00:02:26.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="336" swimtime="00:01:23.59" resultid="8829" heatid="10841" lane="5" entrytime="00:01:23.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="321" swimtime="00:03:01.05" resultid="8830" heatid="10896" lane="3" entrytime="00:03:01.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                    <SPLIT distance="100" swimtime="00:01:28.36" />
                    <SPLIT distance="150" swimtime="00:02:14.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="271" swimtime="00:06:05.18" resultid="8831" heatid="10933" lane="8" entrytime="00:06:10.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                    <SPLIT distance="100" swimtime="00:01:28.21" />
                    <SPLIT distance="150" swimtime="00:02:15.07" />
                    <SPLIT distance="200" swimtime="00:03:01.92" />
                    <SPLIT distance="250" swimtime="00:03:48.39" />
                    <SPLIT distance="300" swimtime="00:04:35.29" />
                    <SPLIT distance="350" swimtime="00:05:21.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-12" firstname="Sasha" gender="M" lastname="Broshevan" nation="POL" athleteid="6109">
              <RESULTS>
                <RESULT eventid="1160" points="412" swimtime="00:00:28.10" resultid="8856" heatid="10708" lane="0" entrytime="00:00:27.00" />
                <RESULT eventid="1190" points="276" swimtime="00:02:55.04" resultid="8857" heatid="10726" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:23.50" />
                    <SPLIT distance="150" swimtime="00:02:15.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="333" swimtime="00:00:34.67" resultid="8858" heatid="10749" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1302" points="410" swimtime="00:01:03.14" resultid="8859" heatid="10785" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="414" swimtime="00:00:30.08" resultid="8860" heatid="10825" lane="5" />
                <RESULT eventid="1452" points="276" swimtime="00:01:19.56" resultid="8861" heatid="10848" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="226" swimtime="00:03:03.50" resultid="8862" heatid="10903" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:01:29.92" />
                    <SPLIT distance="150" swimtime="00:02:18.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="349" swimtime="00:00:37.50" resultid="8863" heatid="10922" lane="1" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Magdalena" gender="F" lastname="Gorostiza" nation="POL" athleteid="6095">
              <RESULTS>
                <RESULT eventid="1287" points="321" swimtime="00:01:15.96" resultid="8845" heatid="10768" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="310" swimtime="00:01:35.01" resultid="8846" heatid="10806" lane="2" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="377" swimtime="00:00:40.79" resultid="8847" heatid="10909" lane="2" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-08" firstname="Przemysław" gender="M" lastname="Osiwała" nation="POL" athleteid="8840">
              <RESULTS>
                <RESULT eventid="1190" points="323" swimtime="00:02:46.04" resultid="8841" heatid="10727" lane="9" entrytime="00:02:40.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:19.37" />
                    <SPLIT distance="150" swimtime="00:02:08.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="296" swimtime="00:02:47.21" resultid="8842" heatid="10795" lane="2" entrytime="00:02:42.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:01:59.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="308" swimtime="00:06:00.91" resultid="8843" heatid="10880" lane="2" entrytime="00:05:38.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:22.76" />
                    <SPLIT distance="150" swimtime="00:02:11.98" />
                    <SPLIT distance="200" swimtime="00:02:59.58" />
                    <SPLIT distance="250" swimtime="00:03:53.21" />
                    <SPLIT distance="300" swimtime="00:04:44.75" />
                    <SPLIT distance="350" swimtime="00:05:23.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="329" swimtime="00:01:12.14" resultid="8844" heatid="10889" lane="5" entrytime="00:01:10.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1347" points="321" swimtime="00:02:35.28" resultid="8866" heatid="10798" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="150" swimtime="00:01:57.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6075" number="1" />
                    <RELAYPOSITION athleteid="6095" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="6108" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="6099" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1497" points="337" swimtime="00:02:18.68" resultid="8867" heatid="10868" lane="8" entrytime="00:02:25.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:06.56" />
                    <SPLIT distance="150" swimtime="00:01:43.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6075" number="1" />
                    <RELAYPOSITION athleteid="6095" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="6099" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="6108" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:03.97" resultid="8864" heatid="10732" lane="2" entrytime="00:02:10.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                    <SPLIT distance="100" swimtime="00:01:01.88" />
                    <SPLIT distance="150" swimtime="00:01:35.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6109" number="1" />
                    <RELAYPOSITION athleteid="6095" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="6075" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="8840" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1653" swimtime="00:02:16.12" resultid="8865" heatid="10928" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:01:21.06" />
                    <SPLIT distance="150" swimtime="00:01:48.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6075" number="1" />
                    <RELAYPOSITION athleteid="6095" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="6081" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="6109" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MALOD" nation="POL" region="05" clubid="4363" name="Masters Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos Rafał" phone="604184311" />
          <ATHLETES>
            <ATHLETE birthdate="1980-04-16" firstname="Joanna" gender="F" lastname="Wilińska-Nowak" nation="POL" athleteid="4387">
              <RESULTS>
                <RESULT eventid="1226" points="360" swimtime="00:00:38.02" resultid="6878" heatid="10738" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1407" points="378" swimtime="00:00:33.77" resultid="6879" heatid="10822" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-11-02" firstname="Ksawery" gender="M" lastname="Wiaderek" nation="POL" athleteid="4392">
              <RESULTS>
                <RESULT eventid="1160" points="501" swimtime="00:00:26.31" resultid="6881" heatid="10707" lane="7" entrytime="00:00:27.00" />
                <RESULT eventid="1242" points="404" swimtime="00:00:32.50" resultid="6882" heatid="10748" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="445" swimtime="00:01:01.42" resultid="6883" heatid="10785" lane="8" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="491" swimtime="00:00:28.42" resultid="6884" heatid="10835" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1578" points="339" swimtime="00:01:11.45" resultid="6885" heatid="10890" lane="7" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-09" firstname="Rafał" gender="M" lastname="Trudnos" nation="POL" athleteid="4381">
              <RESULTS>
                <RESULT eventid="1160" points="415" swimtime="00:00:28.02" resultid="6873" heatid="10705" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1272" points="421" swimtime="00:02:49.40" resultid="6874" heatid="10763" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:19.60" />
                    <SPLIT distance="150" swimtime="00:02:03.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="415" swimtime="00:01:16.54" resultid="6875" heatid="10818" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="394" swimtime="00:00:30.58" resultid="6876" heatid="10834" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1638" points="477" swimtime="00:00:33.80" resultid="6877" heatid="10924" lane="5" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-02" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" athleteid="4412">
              <RESULTS>
                <RESULT eventid="1160" points="448" swimtime="00:00:27.31" resultid="6898" heatid="10709" lane="8" entrytime="00:00:26.00" />
                <RESULT eventid="1302" points="387" swimtime="00:01:04.33" resultid="6899" heatid="10781" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="367" swimtime="00:00:31.32" resultid="6900" heatid="10832" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1638" points="408" swimtime="00:00:35.61" resultid="6901" heatid="10922" lane="2" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-06-12" firstname="Igor" gender="M" lastname="Olejarczyk" nation="POL" athleteid="4375">
              <RESULTS>
                <RESULT eventid="1160" points="454" swimtime="00:00:27.20" resultid="6868" heatid="10706" lane="9" entrytime="00:00:27.50" />
                <RESULT eventid="1332" points="260" swimtime="00:02:54.57" resultid="6869" heatid="10795" lane="6" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:14.43" />
                    <SPLIT distance="150" swimtime="00:02:02.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="436" swimtime="00:00:29.56" resultid="6870" heatid="10836" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1482" points="332" swimtime="00:02:27.28" resultid="6871" heatid="10863" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:09.28" />
                    <SPLIT distance="150" swimtime="00:01:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="397" swimtime="00:01:07.74" resultid="6872" heatid="10890" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-28" firstname="Artur" gender="M" lastname="Frąckowiak" nation="POL" athleteid="4398">
              <RESULTS>
                <RESULT eventid="1128" points="321" swimtime="00:21:11.61" resultid="6886" heatid="10679" lane="7" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:01:56.49" />
                    <SPLIT distance="200" swimtime="00:02:37.00" />
                    <SPLIT distance="250" swimtime="00:03:17.95" />
                    <SPLIT distance="300" swimtime="00:03:58.97" />
                    <SPLIT distance="350" swimtime="00:04:40.00" />
                    <SPLIT distance="400" swimtime="00:05:21.17" />
                    <SPLIT distance="450" swimtime="00:06:02.96" />
                    <SPLIT distance="500" swimtime="00:06:44.66" />
                    <SPLIT distance="550" swimtime="00:07:26.61" />
                    <SPLIT distance="600" swimtime="00:08:08.54" />
                    <SPLIT distance="650" swimtime="00:08:50.81" />
                    <SPLIT distance="700" swimtime="00:09:33.04" />
                    <SPLIT distance="750" swimtime="00:10:16.08" />
                    <SPLIT distance="800" swimtime="00:10:59.17" />
                    <SPLIT distance="850" swimtime="00:11:42.79" />
                    <SPLIT distance="900" swimtime="00:12:26.44" />
                    <SPLIT distance="950" swimtime="00:13:10.02" />
                    <SPLIT distance="1000" swimtime="00:13:53.70" />
                    <SPLIT distance="1050" swimtime="00:14:37.83" />
                    <SPLIT distance="1100" swimtime="00:15:21.81" />
                    <SPLIT distance="1150" swimtime="00:16:06.41" />
                    <SPLIT distance="1200" swimtime="00:16:50.29" />
                    <SPLIT distance="1250" swimtime="00:17:34.52" />
                    <SPLIT distance="1300" swimtime="00:18:18.74" />
                    <SPLIT distance="1350" swimtime="00:19:03.15" />
                    <SPLIT distance="1400" swimtime="00:19:47.24" />
                    <SPLIT distance="1450" swimtime="00:20:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="393" swimtime="00:02:35.53" resultid="6887" heatid="10728" lane="3" entrytime="00:02:33.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:13.16" />
                    <SPLIT distance="150" swimtime="00:02:00.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="463" swimtime="00:01:00.62" resultid="6888" heatid="10784" lane="3" entrytime="00:01:00.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="437" swimtime="00:00:29.55" resultid="6889" heatid="10829" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1482" points="398" swimtime="00:02:18.65" resultid="6890" heatid="10863" lane="2" entrytime="00:02:19.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="100" swimtime="00:01:06.95" />
                    <SPLIT distance="150" swimtime="00:01:43.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="378" swimtime="00:05:04.24" resultid="6891" heatid="10942" lane="6" entrytime="00:05:11.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:11.22" />
                    <SPLIT distance="150" swimtime="00:01:49.35" />
                    <SPLIT distance="200" swimtime="00:02:28.66" />
                    <SPLIT distance="250" swimtime="00:03:07.90" />
                    <SPLIT distance="300" swimtime="00:03:47.45" />
                    <SPLIT distance="350" swimtime="00:04:27.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="4427">
              <RESULTS>
                <RESULT eventid="1098" points="186" swimtime="00:13:11.45" resultid="6910" heatid="10670" lane="5" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:20.10" />
                    <SPLIT distance="150" swimtime="00:02:07.15" />
                    <SPLIT distance="200" swimtime="00:02:57.02" />
                    <SPLIT distance="250" swimtime="00:03:47.26" />
                    <SPLIT distance="300" swimtime="00:04:38.07" />
                    <SPLIT distance="350" swimtime="00:05:30.21" />
                    <SPLIT distance="400" swimtime="00:06:22.16" />
                    <SPLIT distance="450" swimtime="00:07:14.51" />
                    <SPLIT distance="500" swimtime="00:08:06.61" />
                    <SPLIT distance="550" swimtime="00:08:59.48" />
                    <SPLIT distance="600" swimtime="00:09:51.33" />
                    <SPLIT distance="650" swimtime="00:10:42.60" />
                    <SPLIT distance="700" swimtime="00:11:34.17" />
                    <SPLIT distance="750" swimtime="00:12:26.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="322" swimtime="00:00:30.50" resultid="6911" heatid="10695" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1190" points="235" swimtime="00:03:04.53" resultid="6912" heatid="10721" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:26.36" />
                    <SPLIT distance="150" swimtime="00:02:20.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="252" swimtime="00:03:20.83" resultid="6913" heatid="10760" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:01:34.46" />
                    <SPLIT distance="150" swimtime="00:02:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="263" swimtime="00:01:29.13" resultid="6914" heatid="10811" lane="4" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="171" swimtime="00:07:18.99" resultid="6916" heatid="10878" lane="8" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:01:33.56" />
                    <SPLIT distance="150" swimtime="00:02:35.38" />
                    <SPLIT distance="200" swimtime="00:03:35.00" />
                    <SPLIT distance="250" swimtime="00:04:37.62" />
                    <SPLIT distance="300" swimtime="00:05:40.32" />
                    <SPLIT distance="350" swimtime="00:06:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="209" swimtime="00:03:08.42" resultid="6917" heatid="10900" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:28.28" />
                    <SPLIT distance="150" swimtime="00:02:20.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="304" swimtime="00:00:39.26" resultid="6918" heatid="10915" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-18" firstname="Konrad" gender="M" lastname="Hasik" nation="POL" athleteid="4405">
              <RESULTS>
                <RESULT eventid="1190" points="472" swimtime="00:02:26.38" resultid="6892" heatid="10728" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="100" swimtime="00:01:07.03" />
                    <SPLIT distance="150" swimtime="00:01:50.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="482" swimtime="00:00:30.65" resultid="6893" heatid="10751" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1332" points="306" swimtime="00:02:45.42" resultid="6894" heatid="10794" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:58.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="483" swimtime="00:01:06.08" resultid="6895" heatid="10850" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="389" swimtime="00:05:33.81" resultid="6896" heatid="10881" lane="3" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:14.67" />
                    <SPLIT distance="150" swimtime="00:01:58.64" />
                    <SPLIT distance="200" swimtime="00:02:41.91" />
                    <SPLIT distance="250" swimtime="00:03:30.21" />
                    <SPLIT distance="300" swimtime="00:04:17.38" />
                    <SPLIT distance="350" swimtime="00:04:56.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="424" swimtime="00:02:28.94" resultid="6897" heatid="10904" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.75" />
                    <SPLIT distance="150" swimtime="00:01:52.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-14" firstname="Anna" gender="F" lastname="Ostrowska" nation="POL" athleteid="4390">
              <RESULTS>
                <RESULT eventid="1144" points="464" swimtime="00:00:30.65" resultid="6880" heatid="10687" lane="3" entrytime="00:00:30.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-11" firstname="Przemysław" gender="M" lastname="Michniewski" nation="POL" athleteid="4417">
              <RESULTS>
                <RESULT eventid="1160" points="448" swimtime="00:00:27.32" resultid="6902" heatid="10701" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1190" points="389" swimtime="00:02:36.06" resultid="6903" heatid="10725" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="100" swimtime="00:01:11.16" />
                    <SPLIT distance="150" swimtime="00:01:58.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="407" swimtime="00:02:51.25" resultid="6904" heatid="10762" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                    <SPLIT distance="150" swimtime="00:02:05.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="401" swimtime="00:01:17.44" resultid="6905" heatid="10816" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="416" swimtime="00:00:30.03" resultid="6906" heatid="10833" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1638" points="443" swimtime="00:00:34.64" resultid="6907" heatid="10923" lane="2" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-10" firstname="Błażej" gender="M" lastname="Dunajczyk" nation="POL" athleteid="4437">
              <RESULTS>
                <RESULT eventid="1160" points="317" swimtime="00:00:30.66" resultid="6919" heatid="10703" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1302" points="319" swimtime="00:01:08.61" resultid="6920" heatid="10781" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="340" swimtime="00:00:32.11" resultid="6921" heatid="10832" lane="7" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" athleteid="4424">
              <RESULTS>
                <RESULT eventid="1128" points="264" swimtime="00:22:36.22" resultid="6908" heatid="10676" lane="5" entrytime="00:24:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                    <SPLIT distance="100" swimtime="00:01:26.25" />
                    <SPLIT distance="150" swimtime="00:02:11.16" />
                    <SPLIT distance="200" swimtime="00:02:56.23" />
                    <SPLIT distance="250" swimtime="00:03:41.15" />
                    <SPLIT distance="300" swimtime="00:04:26.81" />
                    <SPLIT distance="350" swimtime="00:05:11.80" />
                    <SPLIT distance="400" swimtime="00:05:57.30" />
                    <SPLIT distance="450" swimtime="00:06:42.75" />
                    <SPLIT distance="500" swimtime="00:07:27.86" />
                    <SPLIT distance="550" swimtime="00:08:13.03" />
                    <SPLIT distance="600" swimtime="00:08:58.59" />
                    <SPLIT distance="650" swimtime="00:09:43.47" />
                    <SPLIT distance="700" swimtime="00:10:29.04" />
                    <SPLIT distance="750" swimtime="00:11:15.03" />
                    <SPLIT distance="800" swimtime="00:12:01.17" />
                    <SPLIT distance="850" swimtime="00:12:47.44" />
                    <SPLIT distance="900" swimtime="00:13:33.74" />
                    <SPLIT distance="950" swimtime="00:14:19.84" />
                    <SPLIT distance="1000" swimtime="00:15:05.96" />
                    <SPLIT distance="1050" swimtime="00:15:51.27" />
                    <SPLIT distance="1100" swimtime="00:16:37.06" />
                    <SPLIT distance="1150" swimtime="00:17:23.11" />
                    <SPLIT distance="1200" swimtime="00:18:09.64" />
                    <SPLIT distance="1250" swimtime="00:18:56.19" />
                    <SPLIT distance="1300" swimtime="00:19:42.80" />
                    <SPLIT distance="1350" swimtime="00:20:28.29" />
                    <SPLIT distance="1400" swimtime="00:21:14.31" />
                    <SPLIT distance="1450" swimtime="00:21:56.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="293" swimtime="00:00:31.46" resultid="6909" heatid="10696" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1368" points="471" swimtime="00:02:00.00" resultid="6923" heatid="10802" lane="0" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:04.52" />
                    <SPLIT distance="150" swimtime="00:01:34.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4405" number="1" />
                    <RELAYPOSITION athleteid="4381" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4375" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4392" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1368" points="384" swimtime="00:02:08.50" resultid="6924" heatid="10801" lane="7" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="100" swimtime="00:01:11.13" />
                    <SPLIT distance="150" swimtime="00:01:40.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4427" number="1" />
                    <RELAYPOSITION athleteid="4417" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4398" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4412" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1518" points="497" swimtime="00:01:47.05" resultid="6925" heatid="10872" lane="7" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                    <SPLIT distance="100" swimtime="00:00:54.42" />
                    <SPLIT distance="150" swimtime="00:01:21.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4398" number="1" />
                    <RELAYPOSITION athleteid="4375" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4412" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4392" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1518" points="399" swimtime="00:01:55.17" resultid="6926" heatid="10871" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                    <SPLIT distance="100" swimtime="00:01:00.47" />
                    <SPLIT distance="150" swimtime="00:01:28.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4437" number="1" />
                    <RELAYPOSITION athleteid="4427" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4381" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4417" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:01:55.00" resultid="6922" heatid="10732" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:00:58.86" />
                    <SPLIT distance="150" swimtime="00:01:28.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4387" number="1" />
                    <RELAYPOSITION athleteid="4375" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4390" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4392" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="UCLUB" nation="EST" clubid="3171" name="Meisterujumise U-Klubi">
          <CONTACT email="a_kristiina@hotmail.com" internet="u-klubi.com" name="Kristiina Arusoo" phone="+37256656831" />
          <ATHLETES>
            <ATHLETE birthdate="1954-08-05" firstname="Ossi Albin" gender="M" lastname="Vallemaa" nation="FIN" athleteid="3177">
              <RESULTS>
                <RESULT eventid="1392" points="184" swimtime="00:01:40.37" resultid="6554" heatid="10812" lane="1" entrytime="00:01:36.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="212" swimtime="00:00:44.30" resultid="6555" heatid="10917" lane="9" entrytime="00:00:41.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ASLES" nation="POL" region="WIE" clubid="3346" name="Miejski Klub Pływacki Astromal Leszno" shortname="Miejski Klub Pływacki Astromal">
          <CONTACT email="krzychutomczyk@o2.pl" name="Tomczyk Krzysztof" phone="723524682" />
          <ATHLETES>
            <ATHLETE birthdate="1989-12-20" firstname="Konrad" gender="M" lastname="Nykiel" nation="POL" athleteid="3347">
              <RESULTS>
                <RESULT eventid="1128" points="399" swimtime="00:19:42.62" resultid="6848" heatid="10679" lane="1" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:09.14" />
                    <SPLIT distance="150" swimtime="00:01:47.04" />
                    <SPLIT distance="200" swimtime="00:02:25.98" />
                    <SPLIT distance="250" swimtime="00:03:05.18" />
                    <SPLIT distance="300" swimtime="00:03:44.98" />
                    <SPLIT distance="350" swimtime="00:04:24.79" />
                    <SPLIT distance="400" swimtime="00:05:05.06" />
                    <SPLIT distance="450" swimtime="00:05:45.11" />
                    <SPLIT distance="500" swimtime="00:06:25.24" />
                    <SPLIT distance="550" swimtime="00:07:05.24" />
                    <SPLIT distance="600" swimtime="00:07:45.83" />
                    <SPLIT distance="650" swimtime="00:08:26.25" />
                    <SPLIT distance="700" swimtime="00:09:06.90" />
                    <SPLIT distance="750" swimtime="00:09:47.41" />
                    <SPLIT distance="800" swimtime="00:10:27.34" />
                    <SPLIT distance="850" swimtime="00:11:07.23" />
                    <SPLIT distance="900" swimtime="00:11:47.88" />
                    <SPLIT distance="950" swimtime="00:12:27.95" />
                    <SPLIT distance="1000" swimtime="00:13:08.69" />
                    <SPLIT distance="1050" swimtime="00:13:49.05" />
                    <SPLIT distance="1100" swimtime="00:14:29.54" />
                    <SPLIT distance="1150" swimtime="00:15:09.31" />
                    <SPLIT distance="1200" swimtime="00:15:49.70" />
                    <SPLIT distance="1250" swimtime="00:16:29.43" />
                    <SPLIT distance="1300" swimtime="00:17:09.32" />
                    <SPLIT distance="1350" swimtime="00:17:49.29" />
                    <SPLIT distance="1400" swimtime="00:18:29.30" />
                    <SPLIT distance="1450" swimtime="00:19:07.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="375" swimtime="00:02:37.97" resultid="6849" heatid="10725" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="150" swimtime="00:02:03.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="486" swimtime="00:00:59.63" resultid="6850" heatid="10786" lane="8" entrytime="00:00:59.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="510" swimtime="00:00:28.07" resultid="6851" heatid="10837" lane="9" entrytime="00:00:28.19" />
                <RESULT eventid="1482" points="437" swimtime="00:02:14.40" resultid="6852" heatid="10864" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="6853" heatid="10890" lane="6" entrytime="00:01:07.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-07-14" firstname="Krzysztof" gender="M" lastname="Tomczyk" nation="POL" athleteid="3354">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="6854" heatid="10707" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="6855" heatid="10725" lane="9" entrytime="00:02:50.00" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="6856" heatid="10762" lane="3" entrytime="00:02:55.00" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="6857" heatid="10818" lane="0" entrytime="00:01:16.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="6858" heatid="10923" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-05-02" firstname="Marcin" gender="M" lastname="Kotlarski" nation="POL" athleteid="3360">
              <RESULTS>
                <RESULT eventid="1160" points="456" swimtime="00:00:27.15" resultid="6859" heatid="10708" lane="4" entrytime="00:00:26.38" />
                <RESULT eventid="1190" points="366" swimtime="00:02:39.28" resultid="6860" heatid="10725" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:15.12" />
                    <SPLIT distance="150" swimtime="00:02:02.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="6861" heatid="10786" lane="0" entrytime="00:00:59.50" />
                <RESULT eventid="1482" points="385" swimtime="00:02:20.14" resultid="6862" heatid="10864" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:06.89" />
                    <SPLIT distance="150" swimtime="00:01:43.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" status="DNS" swimtime="00:00:00.00" resultid="6863" heatid="10878" lane="4" entrytime="00:06:30.00" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="6864" heatid="10941" lane="7" entrytime="00:05:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00308" nation="POL" region="08" clubid="2851" name="Mkp Bobry Dębica">
          <CONTACT name="GOGACZ" phone="506694816" />
          <ATHLETES>
            <ATHLETE birthdate="1967-11-09" firstname="Elżbieta" gender="F" lastname="Nowak-Bereś" nation="POL" license="500308600162" athleteid="2869">
              <RESULTS>
                <RESULT eventid="1144" points="155" swimtime="00:00:44.14" resultid="6409" heatid="10682" lane="7" entrytime="00:00:43.50" />
                <RESULT comment="K 14 - Praca nóg  w płaszczyźnie pionowej w dół /z wyjątkiem jednego ruchu po starcie i nawrocie/" eventid="1175" status="DSQ" swimtime="00:04:04.68" resultid="6410" heatid="10713" lane="2" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.79" />
                    <SPLIT distance="100" swimtime="00:02:00.07" />
                    <SPLIT distance="150" swimtime="00:03:10.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="146" swimtime="00:01:38.66" resultid="6411" heatid="10766" lane="2" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="133" swimtime="00:00:47.80" resultid="6412" heatid="10821" lane="8" entrytime="00:00:50.56" />
                <RESULT eventid="1467" points="143" swimtime="00:03:35.96" resultid="6413" heatid="10852" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.81" />
                    <SPLIT distance="100" swimtime="00:01:42.05" />
                    <SPLIT distance="150" swimtime="00:02:39.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="181" swimtime="00:00:52.10" resultid="6414" heatid="10906" lane="3" entrytime="00:00:56.40" />
                <RESULT eventid="1674" points="133" swimtime="00:07:42.72" resultid="6415" heatid="10932" lane="0" entrytime="00:07:34.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.46" />
                    <SPLIT distance="100" swimtime="00:01:45.86" />
                    <SPLIT distance="150" swimtime="00:02:45.55" />
                    <SPLIT distance="200" swimtime="00:03:46.46" />
                    <SPLIT distance="250" swimtime="00:04:47.30" />
                    <SPLIT distance="300" swimtime="00:05:48.08" />
                    <SPLIT distance="350" swimtime="00:06:46.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-11" firstname="Przemysław" gender="M" lastname="Jurek" nation="POL" athleteid="2852">
              <RESULTS>
                <RESULT eventid="1160" points="503" swimtime="00:00:26.28" resultid="6395" heatid="10710" lane="7" entrytime="00:00:25.32" />
                <RESULT eventid="1302" points="516" swimtime="00:00:58.45" resultid="6396" heatid="10787" lane="3" entrytime="00:00:55.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="489" swimtime="00:00:28.47" resultid="6397" heatid="10836" lane="6" entrytime="00:00:28.37" />
                <RESULT eventid="1482" points="459" swimtime="00:02:12.19" resultid="6398" heatid="10866" lane="7" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="100" swimtime="00:01:05.13" />
                    <SPLIT distance="150" swimtime="00:01:39.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="473" swimtime="00:01:03.92" resultid="6399" heatid="10892" lane="9" entrytime="00:01:00.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-07-08" firstname="Andrzej" gender="M" lastname="Maciejczak" nation="POL" athleteid="2862">
              <RESULTS>
                <RESULT eventid="1128" points="181" swimtime="00:25:38.16" resultid="6403" heatid="10675" lane="4" entrytime="00:25:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="100" swimtime="00:01:28.76" />
                    <SPLIT distance="150" swimtime="00:02:20.03" />
                    <SPLIT distance="200" swimtime="00:03:11.68" />
                    <SPLIT distance="250" swimtime="00:04:03.67" />
                    <SPLIT distance="300" swimtime="00:04:55.87" />
                    <SPLIT distance="350" swimtime="00:05:47.28" />
                    <SPLIT distance="400" swimtime="00:06:40.34" />
                    <SPLIT distance="450" swimtime="00:07:31.91" />
                    <SPLIT distance="500" swimtime="00:08:24.48" />
                    <SPLIT distance="550" swimtime="00:09:14.33" />
                    <SPLIT distance="600" swimtime="00:10:06.11" />
                    <SPLIT distance="650" swimtime="00:10:57.66" />
                    <SPLIT distance="700" swimtime="00:11:49.50" />
                    <SPLIT distance="750" swimtime="00:12:40.91" />
                    <SPLIT distance="800" swimtime="00:13:32.90" />
                    <SPLIT distance="850" swimtime="00:14:24.13" />
                    <SPLIT distance="900" swimtime="00:15:16.19" />
                    <SPLIT distance="950" swimtime="00:16:07.19" />
                    <SPLIT distance="1000" swimtime="00:16:59.15" />
                    <SPLIT distance="1050" swimtime="00:17:51.13" />
                    <SPLIT distance="1100" swimtime="00:18:44.00" />
                    <SPLIT distance="1150" swimtime="00:19:35.65" />
                    <SPLIT distance="1200" swimtime="00:20:28.22" />
                    <SPLIT distance="1250" swimtime="00:21:14.07" />
                    <SPLIT distance="1300" swimtime="00:22:13.56" />
                    <SPLIT distance="1350" swimtime="00:23:05.52" />
                    <SPLIT distance="1400" swimtime="00:23:58.40" />
                    <SPLIT distance="1450" swimtime="00:24:49.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="130" swimtime="00:03:44.61" resultid="6404" heatid="10720" lane="5" entrytime="00:03:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:49.10" />
                    <SPLIT distance="150" swimtime="00:03:00.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="196" swimtime="00:01:20.65" resultid="6405" heatid="10776" lane="7" entrytime="00:01:19.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="186" swimtime="00:02:58.62" resultid="6406" heatid="10859" lane="9" entrytime="00:02:56.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="100" swimtime="00:01:24.12" />
                    <SPLIT distance="150" swimtime="00:02:11.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="118" swimtime="00:08:16.39" resultid="6407" heatid="10876" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.26" />
                    <SPLIT distance="100" swimtime="00:02:04.79" />
                    <SPLIT distance="150" swimtime="00:03:12.98" />
                    <SPLIT distance="200" swimtime="00:04:21.62" />
                    <SPLIT distance="250" swimtime="00:05:34.26" />
                    <SPLIT distance="300" swimtime="00:06:42.87" />
                    <SPLIT distance="350" swimtime="00:07:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="185" swimtime="00:06:25.53" resultid="6408" heatid="10938" lane="5" entrytime="00:06:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:01:27.45" />
                    <SPLIT distance="150" swimtime="00:02:16.33" />
                    <SPLIT distance="200" swimtime="00:03:06.57" />
                    <SPLIT distance="250" swimtime="00:03:56.97" />
                    <SPLIT distance="300" swimtime="00:04:47.28" />
                    <SPLIT distance="350" swimtime="00:05:37.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-28" firstname="Sebastian" gender="M" lastname="Gogacz" nation="POL" athleteid="2858">
              <RESULTS>
                <RESULT eventid="1128" points="355" swimtime="00:20:29.68" resultid="6400" heatid="10679" lane="8" entrytime="00:20:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:16.36" />
                    <SPLIT distance="150" swimtime="00:01:57.05" />
                    <SPLIT distance="200" swimtime="00:02:37.74" />
                    <SPLIT distance="250" swimtime="00:03:19.01" />
                    <SPLIT distance="300" swimtime="00:03:59.71" />
                    <SPLIT distance="350" swimtime="00:04:40.63" />
                    <SPLIT distance="400" swimtime="00:05:21.76" />
                    <SPLIT distance="450" swimtime="00:06:02.86" />
                    <SPLIT distance="500" swimtime="00:06:43.07" />
                    <SPLIT distance="550" swimtime="00:07:24.58" />
                    <SPLIT distance="600" swimtime="00:08:04.74" />
                    <SPLIT distance="650" swimtime="00:08:46.04" />
                    <SPLIT distance="700" swimtime="00:09:26.97" />
                    <SPLIT distance="750" swimtime="00:10:07.84" />
                    <SPLIT distance="800" swimtime="00:10:49.06" />
                    <SPLIT distance="850" swimtime="00:11:30.23" />
                    <SPLIT distance="900" swimtime="00:12:11.65" />
                    <SPLIT distance="950" swimtime="00:12:53.14" />
                    <SPLIT distance="1000" swimtime="00:13:34.17" />
                    <SPLIT distance="1050" swimtime="00:14:15.84" />
                    <SPLIT distance="1100" swimtime="00:14:56.76" />
                    <SPLIT distance="1150" swimtime="00:15:38.31" />
                    <SPLIT distance="1200" swimtime="00:16:19.69" />
                    <SPLIT distance="1250" swimtime="00:17:01.93" />
                    <SPLIT distance="1300" swimtime="00:17:43.14" />
                    <SPLIT distance="1350" swimtime="00:18:25.48" />
                    <SPLIT distance="1400" swimtime="00:19:07.30" />
                    <SPLIT distance="1450" swimtime="00:19:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="349" swimtime="00:02:38.31" resultid="6401" heatid="10795" lane="7" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:01:56.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="312" swimtime="00:05:59.43" resultid="6402" heatid="10879" lane="7" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:16.72" />
                    <SPLIT distance="150" swimtime="00:02:06.38" />
                    <SPLIT distance="200" swimtime="00:02:55.92" />
                    <SPLIT distance="250" swimtime="00:03:46.98" />
                    <SPLIT distance="300" swimtime="00:04:39.34" />
                    <SPLIT distance="350" swimtime="00:05:20.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKSZC" nation="POL" region="ZAC" clubid="4606" name="MKP Szczecin">
          <CONTACT email="windmuhle@wp.pl" name="Kowalczyk Piotr" phone="509758055" />
          <ATHLETES>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" athleteid="4627">
              <RESULTS>
                <RESULT eventid="1226" points="256" swimtime="00:00:42.58" resultid="9112" heatid="10736" lane="5" entrytime="00:00:42.70" />
                <RESULT eventid="1437" points="263" swimtime="00:01:30.71" resultid="9113" heatid="10840" lane="3" entrytime="00:01:32.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="255" swimtime="00:03:15.56" resultid="9114" heatid="10896" lane="0" entrytime="00:03:18.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:34.13" />
                    <SPLIT distance="150" swimtime="00:02:24.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="4637">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat F 50-54 lat, międzyczasy na 200dow i 400 dow lepsze od Rekordów Polski Masters w kat. F 50-54 lata" eventid="1059" points="388" swimtime="00:11:04.31" resultid="9120" heatid="10667" lane="5" entrytime="00:10:55.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:16.92" />
                    <SPLIT distance="150" swimtime="00:01:57.79" />
                    <SPLIT distance="200" swimtime="00:02:39.22" />
                    <SPLIT distance="250" swimtime="00:03:20.56" />
                    <SPLIT distance="300" swimtime="00:04:02.13" />
                    <SPLIT distance="350" swimtime="00:04:43.94" />
                    <SPLIT distance="400" swimtime="00:05:26.21" />
                    <SPLIT distance="450" swimtime="00:06:08.34" />
                    <SPLIT distance="500" swimtime="00:06:50.72" />
                    <SPLIT distance="550" swimtime="00:07:33.42" />
                    <SPLIT distance="600" swimtime="00:08:16.08" />
                    <SPLIT distance="650" swimtime="00:08:58.67" />
                    <SPLIT distance="700" swimtime="00:09:41.38" />
                    <SPLIT distance="750" swimtime="00:10:23.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="385" swimtime="00:01:11.52" resultid="9121" heatid="10770" lane="1" entrytime="00:01:10.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat F  50-54  lata" eventid="1467" points="410" swimtime="00:02:32.01" resultid="9122" heatid="10855" lane="8" entrytime="00:02:28.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:13.71" />
                    <SPLIT distance="150" swimtime="00:01:53.12" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1593" points="324" swimtime="00:03:00.47" resultid="9123" heatid="10896" lane="5" entrytime="00:02:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                    <SPLIT distance="100" swimtime="00:01:29.18" />
                    <SPLIT distance="150" swimtime="00:02:15.69" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1674" points="376" swimtime="00:05:27.35" resultid="9124" heatid="10934" lane="1" entrytime="00:05:22.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:17.43" />
                    <SPLIT distance="150" swimtime="00:01:36.44" />
                    <SPLIT distance="250" swimtime="00:01:59.05" />
                    <SPLIT distance="300" swimtime="00:04:04.84" />
                    <SPLIT distance="350" swimtime="00:04:17.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-12" firstname="Zbigniew" gender="M" lastname="Szozda" nation="POL" athleteid="4620">
              <RESULTS>
                <RESULT eventid="1242" points="224" swimtime="00:00:39.54" resultid="9106" heatid="10746" lane="9" entrytime="00:00:38.50" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="9107" heatid="10760" lane="9" entrytime="00:03:26.00" />
                <RESULT eventid="1392" points="238" swimtime="00:01:32.18" resultid="9108" heatid="10814" lane="1" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="199" swimtime="00:01:28.75" resultid="9109" heatid="10847" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="9110" heatid="10887" lane="8" entrytime="00:01:29.00" />
                <RESULT eventid="1638" points="267" swimtime="00:00:41.01" resultid="9111" heatid="10916" lane="5" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-27" firstname="Szymon" gender="M" lastname="Kluczyk" nation="POL" athleteid="4615">
              <RESULTS>
                <RESULT eventid="1098" points="440" swimtime="00:09:54.19" resultid="9102" heatid="10673" lane="2" entrytime="00:09:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:05.68" />
                    <SPLIT distance="150" swimtime="00:01:41.08" />
                    <SPLIT distance="200" swimtime="00:02:17.04" />
                    <SPLIT distance="250" swimtime="00:02:53.52" />
                    <SPLIT distance="300" swimtime="00:03:30.47" />
                    <SPLIT distance="350" swimtime="00:04:07.72" />
                    <SPLIT distance="400" swimtime="00:04:45.41" />
                    <SPLIT distance="450" swimtime="00:05:23.63" />
                    <SPLIT distance="500" swimtime="00:06:02.06" />
                    <SPLIT distance="550" swimtime="00:06:41.32" />
                    <SPLIT distance="600" swimtime="00:07:20.20" />
                    <SPLIT distance="650" swimtime="00:07:59.44" />
                    <SPLIT distance="700" swimtime="00:08:37.53" />
                    <SPLIT distance="750" swimtime="00:09:16.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="334" swimtime="00:02:40.62" resultid="9103" heatid="10795" lane="3" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="100" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:01:56.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="419" swimtime="00:05:25.74" resultid="9104" heatid="10881" lane="9" entrytime="00:05:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:55.64" />
                    <SPLIT distance="200" swimtime="00:02:37.25" />
                    <SPLIT distance="250" swimtime="00:03:25.31" />
                    <SPLIT distance="300" swimtime="00:04:13.91" />
                    <SPLIT distance="350" swimtime="00:04:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="477" swimtime="00:04:41.56" resultid="9105" heatid="10936" lane="8" entrytime="00:10:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-08-21" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="4647">
              <RESULTS>
                <RESULT eventid="1257" points="93" swimtime="00:05:06.51" resultid="9128" heatid="10753" lane="8" entrytime="00:05:06.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.52" />
                    <SPLIT distance="100" swimtime="00:02:31.30" />
                    <SPLIT distance="150" swimtime="00:03:49.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="87" swimtime="00:02:25.16" resultid="9129" heatid="10803" lane="3" entrytime="00:02:30.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="75" swimtime="00:01:09.85" resultid="9130" heatid="10906" lane="9" entrytime="00:01:08.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="4643">
              <RESULTS>
                <RESULT eventid="1272" points="188" swimtime="00:03:41.35" resultid="9125" heatid="10759" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                    <SPLIT distance="100" swimtime="00:01:44.67" />
                    <SPLIT distance="150" swimtime="00:02:42.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="191" swimtime="00:01:39.16" resultid="9126" heatid="10812" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="256" swimtime="00:00:41.59" resultid="9127" heatid="10918" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-02-06" firstname="Lech" gender="M" lastname="Orecki" nation="POL" athleteid="4631">
              <RESULTS>
                <RESULT eventid="1128" points="258" swimtime="00:22:47.05" resultid="9115" heatid="10677" lane="6" entrytime="00:22:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:24.40" />
                    <SPLIT distance="150" swimtime="00:02:10.66" />
                    <SPLIT distance="200" swimtime="00:02:57.80" />
                    <SPLIT distance="250" swimtime="00:03:43.92" />
                    <SPLIT distance="300" swimtime="00:04:30.75" />
                    <SPLIT distance="350" swimtime="00:05:17.47" />
                    <SPLIT distance="400" swimtime="00:06:03.85" />
                    <SPLIT distance="450" swimtime="00:06:50.87" />
                    <SPLIT distance="500" swimtime="00:07:38.55" />
                    <SPLIT distance="550" swimtime="00:08:23.74" />
                    <SPLIT distance="600" swimtime="00:09:09.94" />
                    <SPLIT distance="650" swimtime="00:09:56.15" />
                    <SPLIT distance="700" swimtime="00:10:40.95" />
                    <SPLIT distance="750" swimtime="00:11:25.94" />
                    <SPLIT distance="800" swimtime="00:12:12.31" />
                    <SPLIT distance="850" swimtime="00:12:58.49" />
                    <SPLIT distance="900" swimtime="00:13:45.27" />
                    <SPLIT distance="950" swimtime="00:14:31.75" />
                    <SPLIT distance="1000" swimtime="00:15:18.04" />
                    <SPLIT distance="1050" swimtime="00:16:04.18" />
                    <SPLIT distance="1100" swimtime="00:16:50.15" />
                    <SPLIT distance="1150" swimtime="00:17:34.99" />
                    <SPLIT distance="1200" swimtime="00:18:20.18" />
                    <SPLIT distance="1250" swimtime="00:19:05.71" />
                    <SPLIT distance="1300" swimtime="00:19:51.46" />
                    <SPLIT distance="1350" swimtime="00:20:36.65" />
                    <SPLIT distance="1400" swimtime="00:21:22.53" />
                    <SPLIT distance="1450" swimtime="00:22:06.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="279" swimtime="00:00:31.99" resultid="9116" heatid="10699" lane="9" entrytime="00:00:31.20" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="9117" heatid="10779" lane="5" entrytime="00:01:09.00" />
                <RESULT eventid="1482" points="290" swimtime="00:02:34.06" resultid="9118" heatid="10861" lane="6" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:55.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="9119" heatid="10941" lane="3" entrytime="00:05:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="4607">
              <RESULTS>
                <RESULT eventid="1098" points="340" swimtime="00:10:47.22" resultid="9095" heatid="10672" lane="2" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:14.34" />
                    <SPLIT distance="150" swimtime="00:01:54.42" />
                    <SPLIT distance="200" swimtime="00:02:34.86" />
                    <SPLIT distance="250" swimtime="00:03:15.05" />
                    <SPLIT distance="300" swimtime="00:03:56.23" />
                    <SPLIT distance="350" swimtime="00:04:37.49" />
                    <SPLIT distance="400" swimtime="00:05:18.45" />
                    <SPLIT distance="450" swimtime="00:06:00.37" />
                    <SPLIT distance="500" swimtime="00:06:42.21" />
                    <SPLIT distance="550" swimtime="00:07:24.14" />
                    <SPLIT distance="600" swimtime="00:08:06.09" />
                    <SPLIT distance="650" swimtime="00:08:47.27" />
                    <SPLIT distance="700" swimtime="00:09:29.24" />
                    <SPLIT distance="750" swimtime="00:10:09.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="279" swimtime="00:00:36.75" resultid="9096" heatid="10746" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1452" points="289" swimtime="00:01:18.39" resultid="9098" heatid="10847" lane="3" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="313" swimtime="00:02:44.77" resultid="9100" heatid="10902" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                    <SPLIT distance="100" swimtime="00:01:21.28" />
                    <SPLIT distance="150" swimtime="00:02:04.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="346" swimtime="00:05:13.19" resultid="9101" heatid="10943" lane="0" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:13.76" />
                    <SPLIT distance="150" swimtime="00:01:53.28" />
                    <SPLIT distance="200" swimtime="00:02:34.18" />
                    <SPLIT distance="250" swimtime="00:03:14.69" />
                    <SPLIT distance="300" swimtime="00:03:55.64" />
                    <SPLIT distance="350" swimtime="00:04:35.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1518" points="296" swimtime="00:02:07.19" resultid="9131" heatid="10870" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                    <SPLIT distance="100" swimtime="00:01:03.69" />
                    <SPLIT distance="150" swimtime="00:01:34.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4615" number="1" />
                    <RELAYPOSITION athleteid="4620" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4631" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4643" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="06414" nation="POL" region="14" clubid="9527" name="MKS Piaseczno">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1979-02-21" firstname="Gabriel" gender="M" lastname="Turczyński" nation="POL" athleteid="9528">
              <RESULTS>
                <RESULT eventid="1160" points="532" swimtime="00:00:25.79" resultid="9529" heatid="10710" lane="1" entrytime="00:00:25.43" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01201" nation="POL" region="DOL" clubid="3151" name="MKS Piast Głogów">
          <CONTACT email="skib0303@wp.pl" name="Skiba Tomasz" />
          <ATHLETES>
            <ATHLETE birthdate="1978-08-07" firstname="Krzysztof" gender="M" lastname="Kozakowski" nation="POL" license="101201700273" athleteid="4910">
              <RESULTS>
                <RESULT eventid="1160" points="437" swimtime="00:00:27.55" resultid="6519" heatid="10706" lane="2" entrytime="00:00:27.50" />
                <RESULT eventid="1242" points="342" swimtime="00:00:34.37" resultid="6520" heatid="10747" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1422" points="477" swimtime="00:00:28.69" resultid="6521" heatid="10835" lane="6" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWACA" nation="POL" clubid="3628" name="MKS Swim Academy Termy Jakuba Osawa" shortname="MKS Swim Academy Termy Jakuba ">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1991-01-01" firstname="Agnieszka" gender="F" lastname="Burdelak" nation="POL" athleteid="3629">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="3630" heatid="10674" lane="5" entrytime="00:22:00.00" />
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="3631" heatid="10717" lane="0" entrytime="00:02:58.00" />
                <RESULT eventid="1257" status="DNS" swimtime="00:00:00.00" resultid="3632" heatid="10756" lane="3" entrytime="00:02:58.00" />
                <RESULT eventid="1317" status="DNS" swimtime="00:00:00.00" resultid="3633" heatid="10790" lane="5" entrytime="00:03:00.00" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="3634" heatid="10855" lane="1" entrytime="00:02:25.00" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="3635" heatid="10875" lane="7" entrytime="00:06:00.00" />
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="3636" heatid="10897" lane="0" entrytime="00:02:50.00" />
                <RESULT eventid="1674" status="DNS" swimtime="00:00:00.00" resultid="3637" heatid="10934" lane="8" entrytime="00:05:23.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02711" nation="POL" region="SLA" clubid="3101" name="MOS Dąbrowa Górnicza">
          <CONTACT name="Waliczek Mariusz" phone="606448210" />
          <ATHLETES>
            <ATHLETE birthdate="1997-10-22" firstname="Anna" gender="F" lastname="Teresko" nation="POL" license="102711600109" athleteid="3106">
              <RESULTS>
                <RESULT eventid="1317" points="480" swimtime="00:02:35.57" resultid="6390" heatid="10789" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:11.84" />
                    <SPLIT distance="150" swimtime="00:01:53.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="597" swimtime="00:02:14.16" resultid="6391" heatid="10855" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="150" swimtime="00:01:39.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="6392" heatid="10875" lane="5" entrytime="00:05:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-21" firstname="Patryk" gender="M" lastname="Droś" nation="POL" license="102711200122" athleteid="3102">
              <RESULTS>
                <RESULT eventid="1272" points="582" swimtime="00:02:32.12" resultid="6387" heatid="10764" lane="4" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:13.04" />
                    <SPLIT distance="150" swimtime="00:01:54.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="581" swimtime="00:01:08.45" resultid="6388" heatid="10819" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="553" swimtime="00:00:27.32" resultid="6389" heatid="10838" lane="9" entrytime="00:00:26.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOOST" nation="POL" region="SWI" clubid="2902" name="MOSiR Ostrowiec Św.">
          <CONTACT name="Różalski Józef" phone="510600865" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" license="licencja501012700001" athleteid="2903">
              <RESULTS>
                <RESULT eventid="1098" points="129" swimtime="00:14:54.34" resultid="7771" heatid="10669" lane="2" entrytime="00:19:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.15" />
                    <SPLIT distance="100" swimtime="00:01:39.85" />
                    <SPLIT distance="150" swimtime="00:02:33.99" />
                    <SPLIT distance="200" swimtime="00:03:30.86" />
                    <SPLIT distance="250" swimtime="00:04:27.89" />
                    <SPLIT distance="300" swimtime="00:05:26.28" />
                    <SPLIT distance="350" swimtime="00:06:24.47" />
                    <SPLIT distance="400" swimtime="00:07:21.83" />
                    <SPLIT distance="450" swimtime="00:08:19.55" />
                    <SPLIT distance="500" swimtime="00:09:17.32" />
                    <SPLIT distance="550" swimtime="00:10:08.80" />
                    <SPLIT distance="600" swimtime="00:11:11.58" />
                    <SPLIT distance="650" swimtime="00:12:07.85" />
                    <SPLIT distance="700" swimtime="00:13:05.08" />
                    <SPLIT distance="750" swimtime="00:14:00.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="247" swimtime="00:00:33.31" resultid="7772" heatid="10694" lane="4" entrytime="00:00:35.20" />
                <RESULT eventid="1190" points="137" swimtime="00:03:40.62" resultid="7773" heatid="10720" lane="3" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.60" />
                    <SPLIT distance="100" swimtime="00:01:48.41" />
                    <SPLIT distance="150" swimtime="00:02:52.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="144" swimtime="00:04:02.08" resultid="7774" heatid="10758" lane="7" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.67" />
                    <SPLIT distance="100" swimtime="00:01:57.54" />
                    <SPLIT distance="150" swimtime="00:03:00.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="213" swimtime="00:01:18.54" resultid="7775" heatid="10775" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="133" swimtime="00:01:51.66" resultid="7776" heatid="10810" lane="4" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="235" swimtime="00:00:36.32" resultid="7777" heatid="10828" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1578" points="118" swimtime="00:01:41.31" resultid="7778" heatid="10886" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="196" swimtime="00:00:45.47" resultid="7779" heatid="10914" lane="6" entrytime="00:00:48.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOSTA" nation="POL" region="PDK" clubid="3018" name="MOTYL -SENIOR MOSiR Stalowa Wola" shortname="MOTYL -SENIOR MOSiR Stalowa Wo">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" state="PDKLO" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1949-08-09" firstname="Włodzimierz" gender="M" lastname="Jarzyna" nation="POL" athleteid="3028">
              <RESULTS>
                <RESULT eventid="1098" points="182" swimtime="00:13:17.01" resultid="8060" heatid="10670" lane="0" entrytime="00:13:36.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                    <SPLIT distance="100" swimtime="00:01:36.73" />
                    <SPLIT distance="150" swimtime="00:02:29.62" />
                    <SPLIT distance="200" swimtime="00:03:22.49" />
                    <SPLIT distance="250" swimtime="00:04:14.51" />
                    <SPLIT distance="300" swimtime="00:05:05.89" />
                    <SPLIT distance="350" swimtime="00:05:57.40" />
                    <SPLIT distance="400" swimtime="00:06:48.03" />
                    <SPLIT distance="450" swimtime="00:07:38.02" />
                    <SPLIT distance="500" swimtime="00:08:27.93" />
                    <SPLIT distance="550" swimtime="00:09:18.09" />
                    <SPLIT distance="600" swimtime="00:10:08.57" />
                    <SPLIT distance="650" swimtime="00:10:57.66" />
                    <SPLIT distance="700" swimtime="00:11:46.64" />
                    <SPLIT distance="750" swimtime="00:12:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="246" swimtime="00:00:33.37" resultid="8061" heatid="10697" lane="0" entrytime="00:00:33.15" />
                <RESULT eventid="1190" points="162" swimtime="00:03:29.08" resultid="8062" heatid="10721" lane="0" entrytime="00:03:31.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.69" />
                    <SPLIT distance="100" swimtime="00:01:42.81" />
                    <SPLIT distance="150" swimtime="00:02:47.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="177" swimtime="00:00:42.76" resultid="8063" heatid="10743" lane="5" entrytime="00:00:43.88" />
                <RESULT eventid="1302" points="223" swimtime="00:01:17.26" resultid="8064" heatid="10775" lane="6" entrytime="00:01:22.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="176" swimtime="00:01:32.50" resultid="8065" heatid="10845" lane="4" entrytime="00:01:33.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="152" swimtime="00:07:36.43" resultid="8066" heatid="10877" lane="7" entrytime="00:07:30.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.89" />
                    <SPLIT distance="100" swimtime="00:01:57.66" />
                    <SPLIT distance="150" swimtime="00:02:57.51" />
                    <SPLIT distance="200" swimtime="00:03:54.90" />
                    <SPLIT distance="250" swimtime="00:04:59.27" />
                    <SPLIT distance="300" swimtime="00:06:03.18" />
                    <SPLIT distance="350" swimtime="00:06:51.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="158" swimtime="00:03:26.96" resultid="8067" heatid="10900" lane="3" entrytime="00:03:30.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.74" />
                    <SPLIT distance="100" swimtime="00:01:43.32" />
                    <SPLIT distance="150" swimtime="00:02:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="176" swimtime="00:06:31.97" resultid="8068" heatid="10938" lane="9" entrytime="00:06:38.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.16" />
                    <SPLIT distance="100" swimtime="00:01:35.64" />
                    <SPLIT distance="150" swimtime="00:02:28.46" />
                    <SPLIT distance="200" swimtime="00:03:20.60" />
                    <SPLIT distance="250" swimtime="00:04:11.49" />
                    <SPLIT distance="300" swimtime="00:05:00.11" />
                    <SPLIT distance="350" swimtime="00:05:48.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="3019">
              <RESULTS>
                <RESULT eventid="1128" points="256" swimtime="00:22:50.80" resultid="8052" heatid="10677" lane="0" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                    <SPLIT distance="150" swimtime="00:02:01.72" />
                    <SPLIT distance="200" swimtime="00:02:46.46" />
                    <SPLIT distance="250" swimtime="00:03:31.43" />
                    <SPLIT distance="300" swimtime="00:04:16.49" />
                    <SPLIT distance="350" swimtime="00:05:01.82" />
                    <SPLIT distance="400" swimtime="00:05:47.20" />
                    <SPLIT distance="450" swimtime="00:06:32.88" />
                    <SPLIT distance="500" swimtime="00:07:19.05" />
                    <SPLIT distance="550" swimtime="00:08:05.54" />
                    <SPLIT distance="600" swimtime="00:08:51.99" />
                    <SPLIT distance="650" swimtime="00:09:38.48" />
                    <SPLIT distance="700" swimtime="00:10:24.97" />
                    <SPLIT distance="750" swimtime="00:11:11.79" />
                    <SPLIT distance="800" swimtime="00:11:58.15" />
                    <SPLIT distance="850" swimtime="00:12:45.02" />
                    <SPLIT distance="900" swimtime="00:13:32.56" />
                    <SPLIT distance="950" swimtime="00:14:19.80" />
                    <SPLIT distance="1000" swimtime="00:15:06.62" />
                    <SPLIT distance="1050" swimtime="00:15:53.38" />
                    <SPLIT distance="1100" swimtime="00:16:40.55" />
                    <SPLIT distance="1150" swimtime="00:17:28.19" />
                    <SPLIT distance="1200" swimtime="00:18:14.63" />
                    <SPLIT distance="1250" swimtime="00:19:00.56" />
                    <SPLIT distance="1300" swimtime="00:19:47.06" />
                    <SPLIT distance="1350" swimtime="00:20:33.53" />
                    <SPLIT distance="1400" swimtime="00:21:19.97" />
                    <SPLIT distance="1450" swimtime="00:22:05.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="8053" heatid="10724" lane="3" entrytime="00:02:53.00" />
                <RESULT eventid="1242" points="368" swimtime="00:00:33.54" resultid="8054" heatid="10745" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1272" points="296" swimtime="00:03:10.42" resultid="8055" heatid="10761" lane="9" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                    <SPLIT distance="100" swimtime="00:01:29.72" />
                    <SPLIT distance="150" swimtime="00:02:19.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="303" swimtime="00:01:25.03" resultid="8056" heatid="10813" lane="1" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="314" swimtime="00:01:16.23" resultid="8057" heatid="10847" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="307" swimtime="00:02:45.85" resultid="8058" heatid="10902" lane="8" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:22.18" />
                    <SPLIT distance="150" swimtime="00:02:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="384" swimtime="00:00:36.32" resultid="8059" heatid="10921" lane="1" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="3046">
              <RESULTS>
                <RESULT eventid="1160" points="452" swimtime="00:00:27.24" resultid="8076" heatid="10708" lane="8" entrytime="00:00:26.99" />
                <RESULT eventid="1190" points="499" swimtime="00:02:23.70" resultid="8077" heatid="10730" lane="1" entrytime="00:02:24.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="100" swimtime="00:01:07.10" />
                    <SPLIT distance="150" swimtime="00:01:49.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="516" swimtime="00:00:58.45" resultid="8078" heatid="10787" lane="1" entrytime="00:00:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="504" swimtime="00:00:28.18" resultid="8079" heatid="10837" lane="1" entrytime="00:00:27.99" />
                <RESULT eventid="1482" points="490" swimtime="00:02:09.35" resultid="8080" heatid="10866" lane="0" entrytime="00:02:07.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                    <SPLIT distance="100" swimtime="00:01:02.81" />
                    <SPLIT distance="150" swimtime="00:01:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="522" swimtime="00:01:01.86" resultid="8081" heatid="10891" lane="4" entrytime="00:01:00.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="497" swimtime="00:04:37.73" resultid="8082" heatid="10945" lane="7" entrytime="00:04:39.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:06.24" />
                    <SPLIT distance="150" swimtime="00:01:41.75" />
                    <SPLIT distance="200" swimtime="00:02:17.36" />
                    <SPLIT distance="250" swimtime="00:02:52.95" />
                    <SPLIT distance="300" swimtime="00:03:28.61" />
                    <SPLIT distance="350" swimtime="00:04:03.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="3038">
              <RESULTS>
                <RESULT eventid="1144" points="294" swimtime="00:00:35.66" resultid="8069" heatid="10684" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1175" points="276" swimtime="00:03:13.51" resultid="8070" heatid="10715" lane="1" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                    <SPLIT distance="100" swimtime="00:01:34.40" />
                    <SPLIT distance="150" swimtime="00:02:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="263" swimtime="00:03:37.06" resultid="8071" heatid="10754" lane="4" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.10" />
                    <SPLIT distance="100" swimtime="00:01:46.27" />
                    <SPLIT distance="150" swimtime="00:02:43.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="269" swimtime="00:00:37.82" resultid="8072" heatid="10822" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="8073" heatid="10874" lane="8" entrytime="00:07:05.00" />
                <RESULT eventid="1562" points="183" swimtime="00:01:37.63" resultid="8074" heatid="10883" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="250" swimtime="00:00:46.75" resultid="8075" heatid="10908" lane="8" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EULVI" nation="UKR" clubid="4951" name="MSC Euro-Lviv">
          <CONTACT city="Lviv" email="riff@mail.lviv.ua" fax="+48 537 723 854" internet="www.mastersswim.com.ua" name="Ruslan FRIAUF" phone="+38 067 673 47 96" zip="79012" />
          <ATHLETES>
            <ATHLETE birthdate="1976-02-03" firstname="Romana" gender="F" lastname="Sirenko" nation="UKR" athleteid="6987">
              <RESULTS>
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="6988" heatid="10715" lane="4" entrytime="00:03:10.00" />
                <RESULT eventid="1226" status="DNS" swimtime="00:00:00.00" resultid="6989" heatid="10737" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="1407" status="DNS" swimtime="00:00:00.00" resultid="6990" heatid="10822" lane="5" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-18" firstname="Dmytro" gender="M" lastname="Melnyk" nation="UKR" athleteid="6967">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="6968" heatid="10707" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="6969" heatid="10784" lane="5" entrytime="00:01:00.50" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="6970" heatid="10817" lane="3" entrytime="00:01:17.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="6971" heatid="10924" lane="7" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-11-03" firstname="Volodymyr" gender="M" lastname="Ivat" nation="UKR" athleteid="6972">
              <RESULTS>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="6973" heatid="10763" lane="9" entrytime="00:02:51.00" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="6974" heatid="10817" lane="5" entrytime="00:01:17.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="6975" heatid="10890" lane="3" entrytime="00:01:07.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="6976" heatid="10924" lane="8" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-18" firstname="Ihor" gender="M" lastname="Shchotkin" nation="UKR" athleteid="6977">
              <RESULTS>
                <RESULT eventid="1160" points="539" swimtime="00:00:25.69" resultid="6978" heatid="10710" lane="2" entrytime="00:00:25.10" />
                <RESULT eventid="1302" points="515" swimtime="00:00:58.49" resultid="6979" heatid="10786" lane="5" entrytime="00:00:58.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="514" swimtime="00:00:27.99" resultid="6980" heatid="10837" lane="3" entrytime="00:00:27.50" />
                <RESULT eventid="1638" points="508" swimtime="00:00:33.10" resultid="6981" heatid="10925" lane="4" entrytime="00:00:31.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-13" firstname="Oleksandr" gender="M" lastname="Syrbu" nation="UKR" athleteid="6982">
              <RESULTS>
                <RESULT eventid="1160" points="478" swimtime="00:00:26.74" resultid="6983" heatid="10708" lane="3" entrytime="00:00:26.50" />
                <RESULT eventid="1332" points="404" swimtime="00:02:30.72" resultid="6984" heatid="10796" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:12.19" />
                    <SPLIT distance="150" swimtime="00:01:51.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="548" swimtime="00:00:27.40" resultid="6985" heatid="10837" lane="7" entrytime="00:00:27.60" />
                <RESULT eventid="1578" points="390" swimtime="00:01:08.18" resultid="6986" heatid="10891" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-13" firstname="Bogdan" gender="M" lastname="Osidach" nation="UKR" athleteid="6965">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="6966" heatid="10699" lane="6" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-03-31" firstname="Myron" gender="M" lastname="Kolodko" nation="UKR" athleteid="6045" />
            <ATHLETE birthdate="1969-01-07" firstname="Ruslan" gender="M" lastname="Friauf" nation="UKR" athleteid="6991">
              <RESULTS>
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="6992" heatid="10745" lane="4" entrytime="00:00:38.60" />
                <RESULT eventid="1452" status="DNS" swimtime="00:00:00.00" resultid="6993" heatid="10846" lane="4" entrytime="00:01:25.50" />
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="6994" heatid="10901" lane="5" entrytime="00:03:05.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00403" nation="POL" region="03" clubid="2827" name="MUKS Lider Chełm">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1941-10-11" firstname="Janusz" gender="M" lastname="Golik" nation="POL" license="100403700118" athleteid="2828">
              <RESULTS>
                <RESULT eventid="1272" points="125" swimtime="00:04:13.82" resultid="6371" heatid="10758" lane="8" entrytime="00:04:10.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.78" />
                    <SPLIT distance="100" swimtime="00:02:08.41" />
                    <SPLIT distance="150" swimtime="00:03:14.75" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn w  kat K  75-79  lat" eventid="1332" points="54" swimtime="00:04:53.58" resultid="6372" heatid="10792" lane="8" entrytime="00:04:53.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.45" />
                    <SPLIT distance="100" swimtime="00:02:23.33" />
                    <SPLIT distance="150" swimtime="00:03:43.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="150" swimtime="00:01:47.45" resultid="6373" heatid="10811" lane="8" entrytime="00:01:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="81" swimtime="00:00:51.68" resultid="6374" heatid="10826" lane="4" entrytime="00:00:47.15" />
                <RESULT eventid="1578" points="72" swimtime="00:01:59.73" resultid="6375" heatid="10886" lane="9" entrytime="00:01:52.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="198" swimtime="00:00:45.29" resultid="6376" heatid="10915" lane="2" entrytime="00:00:45.09" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06611" nation="POL" region="SLA" clubid="6036" name="Młodzieżowy Klub Pływacki Wodnik 29 Tychy" shortname="Młodzieżowy Klub Pływacki Wodn">
          <CONTACT city="Tychy" email="marekmrozw29@gmail.com" internet="www.wodnik29.pl" name="Marek Mróz" phone="782985239" state="SLA" street="Damrota 170" zip="43-100" />
          <ATHLETES>
            <ATHLETE birthdate="1995-07-13" firstname="Szymon" gender="M" lastname="Warwas" nation="POL" athleteid="6037">
              <RESULTS>
                <RESULT eventid="1160" points="614" swimtime="00:00:24.60" resultid="8415" heatid="10711" lane="6" entrytime="00:00:24.40" />
                <RESULT eventid="1242" points="527" swimtime="00:00:29.75" resultid="8416" heatid="10751" lane="4" entrytime="00:00:27.80" />
                <RESULT eventid="1302" points="590" swimtime="00:00:55.91" resultid="8417" heatid="10787" lane="4" entrytime="00:00:55.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="618" swimtime="00:00:26.32" resultid="8418" heatid="10838" lane="2" entrytime="00:00:25.80" />
                <RESULT eventid="1452" points="464" swimtime="00:01:06.93" resultid="8419" heatid="10850" lane="5" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="464" swimtime="00:01:04.35" resultid="8420" heatid="10892" lane="3" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="420" swimtime="00:00:35.26" resultid="8421" heatid="10923" lane="4" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NADEC" nation="POL" region="14" clubid="4982" name="Nabaiji Team Decathlon">
          <CONTACT city="Toruń" email="filip.wojciechowski@decathlon.com" name="Filip Wojciechowski" phone="503414875" state="KP" street="Żółkiewskiego 15" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1987-05-17" firstname="Zuzanna" gender="F" lastname="Kacalska" nation="POL" athleteid="4983">
              <RESULTS>
                <RESULT eventid="1144" points="401" swimtime="00:00:32.16" resultid="7078" heatid="10686" lane="5" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1287" points="398" swimtime="00:01:10.77" resultid="7079" heatid="10769" lane="3" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="403" swimtime="00:02:32.88" resultid="7080" heatid="10854" lane="5" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:13.35" />
                    <SPLIT distance="150" swimtime="00:01:53.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-02-20" firstname="Maciej" gender="M" lastname="Jekiełek" nation="POL" athleteid="4996">
              <RESULTS>
                <RESULT eventid="1160" points="465" swimtime="00:00:26.98" resultid="7089" heatid="10709" lane="7" entrytime="00:00:26.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-04-06" firstname="Martyna" gender="F" lastname="Górajewska" nation="POL" athleteid="4998">
              <RESULTS>
                <RESULT eventid="1376" points="366" swimtime="00:01:29.94" resultid="7090" heatid="10807" lane="4" entrytime="00:01:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="369" swimtime="00:00:41.08" resultid="7091" heatid="10910" lane="7" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1144" points="418" swimtime="00:00:31.72" resultid="9374" heatid="10687" lane="6" entrytime="00:00:30.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-06" firstname="Paweł" gender="M" lastname="Bednarczyk" nation="POL" athleteid="4987">
              <RESULTS>
                <RESULT eventid="1160" points="644" swimtime="00:00:24.21" resultid="7081" heatid="10710" lane="3" entrytime="00:00:25.00" entrycourse="LCM" />
                <RESULT eventid="1190" points="495" swimtime="00:02:24.04" resultid="7082" heatid="10730" lane="2" entrytime="00:02:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                    <SPLIT distance="100" swimtime="00:01:07.69" />
                    <SPLIT distance="150" swimtime="00:01:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="638" swimtime="00:00:54.48" resultid="7083" heatid="10788" lane="2" entrytime="00:00:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="387" swimtime="00:02:32.96" resultid="7084" heatid="10796" lane="1" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:11.83" />
                    <SPLIT distance="150" swimtime="00:01:51.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="660" swimtime="00:00:25.76" resultid="7085" heatid="10838" lane="5" entrytime="00:00:25.50" entrycourse="LCM" />
                <RESULT eventid="1482" points="501" swimtime="00:02:08.35" resultid="7086" heatid="10865" lane="4" entrytime="00:02:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                    <SPLIT distance="100" swimtime="00:01:01.31" />
                    <SPLIT distance="150" swimtime="00:01:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="624" swimtime="00:00:58.29" resultid="7087" heatid="10892" lane="8" entrytime="00:01:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="451" swimtime="00:04:46.91" resultid="7088" heatid="10935" lane="7" entrytime="00:04:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:06.07" />
                    <SPLIT distance="150" swimtime="00:01:41.93" />
                    <SPLIT distance="200" swimtime="00:02:19.23" />
                    <SPLIT distance="250" swimtime="00:02:56.34" />
                    <SPLIT distance="300" swimtime="00:03:34.20" />
                    <SPLIT distance="350" swimtime="00:04:11.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-20" firstname="Rafał" gender="M" lastname="Liszewski" nation="POL" athleteid="5001">
              <RESULTS>
                <RESULT eventid="1160" points="444" swimtime="00:00:27.40" resultid="7092" heatid="10707" lane="4" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="1242" points="403" swimtime="00:00:32.52" resultid="7093" heatid="10749" lane="3" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="7094" heatid="10834" lane="4" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1638" points="552" swimtime="00:00:32.19" resultid="7095" heatid="10924" lane="1" entrytime="00:00:34.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" status="EXH" swimtime="00:01:55.88" resultid="7096" heatid="10731" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                    <SPLIT distance="100" swimtime="00:00:58.56" />
                    <SPLIT distance="150" swimtime="00:01:30.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4996" number="1" />
                    <RELAYPOSITION athleteid="4998" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4983" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4987" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1653" swimtime="00:02:13.09" resultid="7097" heatid="10927" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="150" swimtime="00:01:41.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5001" number="1" />
                    <RELAYPOSITION athleteid="4998" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4987" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4983" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NEPRA" nation="CZE" clubid="3638" name="Neptun Masters Praha">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1968-01-01" firstname="Hana" gender="F" lastname="Bohuslávková" nation="CZE" athleteid="3645">
              <RESULTS>
                <RESULT eventid="1175" points="400" swimtime="00:02:51.10" resultid="3646" heatid="10717" lane="1" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:19.08" />
                    <SPLIT distance="150" swimtime="00:02:08.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="450" swimtime="00:03:01.46" resultid="3647" heatid="10756" lane="7" entrytime="00:03:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:01:27.41" />
                    <SPLIT distance="150" swimtime="00:02:13.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="473" swimtime="00:01:22.55" resultid="3648" heatid="10808" lane="5" entrytime="00:01:22.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="457" swimtime="00:00:38.25" resultid="3649" heatid="10911" lane="8" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Tomáš" gender="M" lastname="Vonšovský" nation="CZE" athleteid="3656">
              <RESULTS>
                <RESULT eventid="1242" points="361" swimtime="00:00:33.75" resultid="3657" heatid="10749" lane="8" entrytime="00:00:32.57" />
                <RESULT eventid="1422" points="406" swimtime="00:00:30.27" resultid="3658" heatid="10834" lane="8" entrytime="00:00:30.38" />
                <RESULT eventid="1578" points="380" swimtime="00:01:08.73" resultid="3659" heatid="10890" lane="2" entrytime="00:01:08.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Denis" gender="M" lastname="Bushkov" nation="CZE" athleteid="3639">
              <RESULTS>
                <RESULT eventid="1098" points="452" swimtime="00:09:49.06" resultid="3640" heatid="10673" lane="1" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:46.57" />
                    <SPLIT distance="200" swimtime="00:02:23.23" />
                    <SPLIT distance="250" swimtime="00:03:00.23" />
                    <SPLIT distance="300" swimtime="00:03:37.53" />
                    <SPLIT distance="350" swimtime="00:04:14.96" />
                    <SPLIT distance="400" swimtime="00:04:52.64" />
                    <SPLIT distance="450" swimtime="00:05:29.67" />
                    <SPLIT distance="500" swimtime="00:06:06.94" />
                    <SPLIT distance="550" swimtime="00:06:44.41" />
                    <SPLIT distance="600" swimtime="00:07:21.93" />
                    <SPLIT distance="650" swimtime="00:07:59.03" />
                    <SPLIT distance="700" swimtime="00:08:36.20" />
                    <SPLIT distance="750" swimtime="00:09:13.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="408" swimtime="00:02:33.68" resultid="3641" heatid="10728" lane="1" entrytime="00:02:35.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="150" swimtime="00:01:58.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="305" swimtime="00:02:45.65" resultid="3642" heatid="10794" lane="2" entrytime="00:02:55.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:17.79" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="463" swimtime="00:02:11.83" resultid="3643" heatid="10864" lane="9" entrytime="00:02:15.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                    <SPLIT distance="100" swimtime="00:01:03.57" />
                    <SPLIT distance="150" swimtime="00:01:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="480" swimtime="00:04:40.90" resultid="3644" heatid="10944" lane="6" entrytime="00:04:50.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:06.80" />
                    <SPLIT distance="150" swimtime="00:01:42.03" />
                    <SPLIT distance="200" swimtime="00:02:17.79" />
                    <SPLIT distance="250" swimtime="00:02:53.60" />
                    <SPLIT distance="300" swimtime="00:03:29.80" />
                    <SPLIT distance="350" swimtime="00:04:05.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Pavla" gender="F" lastname="Duplinska" nation="CZE" athleteid="3650">
              <RESULTS>
                <RESULT eventid="1144" points="86" swimtime="00:00:53.75" resultid="3651" heatid="10681" lane="3" entrytime="00:00:55.03" />
                <RESULT eventid="1226" points="95" swimtime="00:00:59.30" resultid="3652" heatid="10735" lane="9" entrytime="00:00:59.75" />
                <RESULT eventid="1287" points="57" swimtime="00:02:14.97" resultid="3653" heatid="10765" lane="4" entrytime="00:02:04.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="51" swimtime="00:01:05.56" resultid="3654" heatid="10820" lane="5" entrytime="00:00:57.80" />
                <RESULT eventid="1437" points="84" swimtime="00:02:12.43" resultid="3655" heatid="10839" lane="2" entrytime="00:02:14.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCNEW" nation="GBR" clubid="9052" name="Newmarket and District SC">
          <ATHLETES>
            <ATHLETE birthdate="1966-01-01" firstname="Lisa" gender="F" lastname="Withers" nation="GBR" athleteid="3791">
              <RESULTS>
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="3792" heatid="10684" lane="3" entrytime="00:00:35.68" />
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="3793" heatid="10716" lane="8" entrytime="00:03:09.43" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIBIAL" nation="BLR" clubid="5816" name="Niezrzeszony">
          <CONTACT name="s" />
          <ATHLETES>
            <ATHLETE birthdate="1950-01-01" firstname="Kuzmina" gender="F" lastname="Nadzeya" nation="BLR" athleteid="5822">
              <RESULTS>
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="7326" heatid="10682" lane="2" entrytime="00:00:43.50" />
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="7327" heatid="10906" lane="1" entrytime="00:01:00.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yury" gender="M" lastname="Komov" nameprefix="a" nation="BLR" athleteid="5817">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="7322" heatid="10694" lane="5" entrytime="00:00:35.20" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="7323" heatid="10759" lane="0" entrytime="00:03:35.50" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="7324" heatid="10812" lane="7" entrytime="00:01:36.50" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="7325" heatid="10917" lane="0" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEZR" nation="POL" region="14" clubid="3379" name="Niezrzeszony">
          <CONTACT name="Błazucka" />
          <ATHLETES>
            <ATHLETE birthdate="1962-01-01" firstname="Michał" gender="M" lastname="Biały" nation="POL" athleteid="10615">
              <RESULTS>
                <RESULT eventid="1190" points="247" swimtime="00:03:01.47" resultid="10616" heatid="10719" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:25.40" />
                    <SPLIT distance="150" swimtime="00:02:17.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="202" swimtime="00:00:40.95" resultid="10617" heatid="10740" lane="7" />
                <RESULT eventid="1452" points="188" swimtime="00:01:30.43" resultid="10618" heatid="10843" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Ireneusz" gender="M" lastname="Stachurski" nation="POL" athleteid="7291">
              <RESULTS>
                <RESULT eventid="1160" points="182" swimtime="00:00:36.89" resultid="9813" heatid="10692" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="9814" heatid="10774" lane="1" entrytime="00:01:30.00" />
                <RESULT eventid="1422" points="88" swimtime="00:00:50.30" resultid="9815" heatid="10826" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="9816" heatid="10858" lane="8" entrytime="00:03:10.00" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="9817" heatid="10937" lane="0" entrytime="00:07:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Bernard" gender="M" lastname="Wierzbik" nation="POL" athleteid="7221">
              <RESULTS>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="10272" heatid="10723" lane="9" entrytime="00:03:07.00" />
                <RESULT eventid="1332" points="190" swimtime="00:03:13.69" resultid="10273" heatid="10793" lane="2" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                    <SPLIT distance="100" swimtime="00:01:28.99" />
                    <SPLIT distance="150" swimtime="00:02:22.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="286" swimtime="00:00:34.03" resultid="10274" heatid="10830" lane="8" entrytime="00:00:34.50" />
                <RESULT eventid="1546" points="225" swimtime="00:06:40.33" resultid="10275" heatid="10878" lane="2" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:01:29.23" />
                    <SPLIT distance="200" swimtime="00:03:17.24" />
                    <SPLIT distance="250" swimtime="00:04:13.14" />
                    <SPLIT distance="300" swimtime="00:05:10.05" />
                    <SPLIT distance="350" swimtime="00:05:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="230" swimtime="00:01:21.25" resultid="10276" heatid="10887" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="Maja" gender="F" lastname="Krzysiek" nation="POL" athleteid="7252">
              <RESULTS>
                <RESULT eventid="1175" points="331" swimtime="00:03:02.29" resultid="10294" heatid="10715" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:01:28.94" />
                    <SPLIT distance="150" swimtime="00:02:17.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="422" swimtime="00:01:25.75" resultid="10295" heatid="10808" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="429" swimtime="00:00:39.07" resultid="10296" heatid="10909" lane="5" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Dymitr" gender="M" lastname="Bielskyi" nation="POL" athleteid="10619">
              <RESULTS>
                <RESULT eventid="1272" points="312" swimtime="00:03:07.08" resultid="10620" heatid="10761" lane="0" entrytime="00:03:10.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                    <SPLIT distance="100" swimtime="00:01:30.39" />
                    <SPLIT distance="150" swimtime="00:02:19.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="315" swimtime="00:01:23.90" resultid="10621" heatid="10815" lane="5" entrytime="00:01:24.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="188" swimtime="00:02:57.86" resultid="10622" heatid="10859" lane="3" entrytime="00:02:50.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                    <SPLIT distance="150" swimtime="00:02:12.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Filip" gender="M" lastname="Gawłowski" nation="POL" athleteid="9790">
              <RESULTS>
                <RESULT eventid="1160" points="138" swimtime="00:00:40.39" resultid="9791" heatid="10691" lane="1" entrytime="00:00:46.50" />
                <RESULT eventid="1392" points="156" swimtime="00:01:45.92" resultid="9792" heatid="10810" lane="2" entrytime="00:01:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="218" swimtime="00:00:43.87" resultid="9793" heatid="10913" lane="5" entrytime="00:00:53.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Sigitas" gender="M" lastname="Katkevicius" nation="POL" athleteid="7317">
              <RESULTS>
                <RESULT eventid="1160" points="356" swimtime="00:00:29.50" resultid="10329" heatid="10701" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1242" points="289" swimtime="00:00:36.33" resultid="10330" heatid="10746" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1392" points="300" swimtime="00:01:25.29" resultid="10331" heatid="10814" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="354" swimtime="00:00:37.32" resultid="10332" heatid="10920" lane="3" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Wawrzyniec" gender="M" lastname="Ambroziak" nation="POL" athleteid="7198">
              <RESULTS>
                <RESULT eventid="1160" points="500" swimtime="00:00:26.33" resultid="9806" heatid="10709" lane="9" entrytime="00:00:26.30" />
                <RESULT eventid="1422" points="502" swimtime="00:00:28.22" resultid="9807" heatid="10836" lane="4" entrytime="00:00:28.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Tomasz" gender="M" lastname="Spychalski" nation="POL" athleteid="9368">
              <RESULTS>
                <RESULT eventid="1128" points="305" swimtime="00:21:32.86" resultid="10640" heatid="10677" lane="4" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:15.70" />
                    <SPLIT distance="150" swimtime="00:01:57.66" />
                    <SPLIT distance="200" swimtime="00:02:40.18" />
                    <SPLIT distance="250" swimtime="00:03:23.29" />
                    <SPLIT distance="300" swimtime="00:04:06.19" />
                    <SPLIT distance="350" swimtime="00:04:48.99" />
                    <SPLIT distance="400" swimtime="00:05:32.94" />
                    <SPLIT distance="450" swimtime="00:06:16.49" />
                    <SPLIT distance="500" swimtime="00:07:00.09" />
                    <SPLIT distance="550" swimtime="00:07:43.93" />
                    <SPLIT distance="600" swimtime="00:08:28.05" />
                    <SPLIT distance="650" swimtime="00:09:11.45" />
                    <SPLIT distance="700" swimtime="00:09:55.37" />
                    <SPLIT distance="750" swimtime="00:10:38.88" />
                    <SPLIT distance="800" swimtime="00:11:23.04" />
                    <SPLIT distance="850" swimtime="00:12:06.43" />
                    <SPLIT distance="900" swimtime="00:12:50.55" />
                    <SPLIT distance="950" swimtime="00:13:34.36" />
                    <SPLIT distance="1000" swimtime="00:14:18.10" />
                    <SPLIT distance="1050" swimtime="00:15:02.04" />
                    <SPLIT distance="1100" swimtime="00:15:46.05" />
                    <SPLIT distance="1150" swimtime="00:16:29.73" />
                    <SPLIT distance="1200" swimtime="00:17:13.98" />
                    <SPLIT distance="1250" swimtime="00:17:57.97" />
                    <SPLIT distance="1300" swimtime="00:18:42.39" />
                    <SPLIT distance="1350" swimtime="00:19:26.58" />
                    <SPLIT distance="1400" swimtime="00:20:11.27" />
                    <SPLIT distance="1450" swimtime="00:20:54.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="David" gender="M" lastname="Kochwasser" nation="POL" athleteid="7164">
              <RESULTS>
                <RESULT eventid="1160" points="367" swimtime="00:00:29.19" resultid="10230" heatid="10702" lane="1" entrytime="00:00:29.25" />
                <RESULT eventid="1302" points="347" swimtime="00:01:06.75" resultid="10231" heatid="10780" lane="7" entrytime="00:01:07.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="294" swimtime="00:01:25.90" resultid="10232" heatid="10815" lane="1" entrytime="00:01:25.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="358" swimtime="00:00:31.56" resultid="10233" heatid="10830" lane="4" entrytime="00:00:33.45" />
                <RESULT eventid="1638" points="364" swimtime="00:00:37.00" resultid="10234" heatid="10920" lane="0" entrytime="00:00:38.63" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Šíp" gender="M" lastname="Jiří" nation="POL" athleteid="10235">
              <RESULTS>
                <RESULT eventid="1160" points="428" swimtime="00:00:27.73" resultid="10236" heatid="10705" lane="5" entrytime="00:00:27.70" />
                <RESULT eventid="1190" points="377" swimtime="00:02:37.76" resultid="10237" heatid="10726" lane="3" entrytime="00:02:41.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:14.64" />
                    <SPLIT distance="150" swimtime="00:02:02.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="382" swimtime="00:00:33.13" resultid="10238" heatid="10749" lane="0" entrytime="00:00:32.90" />
                <RESULT eventid="1302" points="470" swimtime="00:01:00.32" resultid="10239" heatid="10784" lane="6" entrytime="00:01:00.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="377" swimtime="00:01:11.72" resultid="10240" heatid="10848" lane="4" entrytime="00:01:11.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="330" swimtime="00:02:41.81" resultid="10241" heatid="10903" lane="8" entrytime="00:02:43.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:17.66" />
                    <SPLIT distance="150" swimtime="00:02:00.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Łukasz" gender="M" lastname="Chmiel" nation="POL" athleteid="7261">
              <RESULTS>
                <RESULT eventid="1098" points="414" swimtime="00:10:06.34" resultid="10302" heatid="10673" lane="4" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:05.82" />
                    <SPLIT distance="150" swimtime="00:01:42.07" />
                    <SPLIT distance="200" swimtime="00:02:19.05" />
                    <SPLIT distance="250" swimtime="00:02:56.46" />
                    <SPLIT distance="300" swimtime="00:03:34.66" />
                    <SPLIT distance="350" swimtime="00:04:13.50" />
                    <SPLIT distance="400" swimtime="00:04:52.88" />
                    <SPLIT distance="450" swimtime="00:05:32.23" />
                    <SPLIT distance="500" swimtime="00:06:12.62" />
                    <SPLIT distance="550" swimtime="00:06:52.45" />
                    <SPLIT distance="600" swimtime="00:07:32.79" />
                    <SPLIT distance="650" swimtime="00:08:13.07" />
                    <SPLIT distance="700" swimtime="00:08:52.81" />
                    <SPLIT distance="750" swimtime="00:09:31.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" status="DSQ" swimtime="00:20:46.59" resultid="10303" heatid="10679" lane="4" entrytime="00:17:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="150" swimtime="00:01:54.07" />
                    <SPLIT distance="200" swimtime="00:02:35.07" />
                    <SPLIT distance="250" swimtime="00:03:15.92" />
                    <SPLIT distance="300" swimtime="00:03:58.10" />
                    <SPLIT distance="350" swimtime="00:04:39.85" />
                    <SPLIT distance="400" swimtime="00:05:21.74" />
                    <SPLIT distance="450" swimtime="00:06:03.89" />
                    <SPLIT distance="500" swimtime="00:06:46.57" />
                    <SPLIT distance="550" swimtime="00:07:29.25" />
                    <SPLIT distance="600" swimtime="00:08:11.40" />
                    <SPLIT distance="650" swimtime="00:08:53.48" />
                    <SPLIT distance="700" swimtime="00:09:35.32" />
                    <SPLIT distance="750" swimtime="00:10:16.89" />
                    <SPLIT distance="800" swimtime="00:10:59.16" />
                    <SPLIT distance="850" swimtime="00:11:41.22" />
                    <SPLIT distance="900" swimtime="00:12:23.22" />
                    <SPLIT distance="950" swimtime="00:13:04.83" />
                    <SPLIT distance="1000" swimtime="00:13:46.66" />
                    <SPLIT distance="1050" swimtime="00:14:28.45" />
                    <SPLIT distance="1100" swimtime="00:15:11.25" />
                    <SPLIT distance="1150" swimtime="00:15:53.61" />
                    <SPLIT distance="1200" swimtime="00:16:36.36" />
                    <SPLIT distance="1250" swimtime="00:17:18.65" />
                    <SPLIT distance="1300" swimtime="00:18:01.96" />
                    <SPLIT distance="1350" swimtime="00:18:36.66" />
                    <SPLIT distance="1400" swimtime="00:19:25.10" />
                    <SPLIT distance="1450" swimtime="00:20:06.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="10304" heatid="10711" lane="1" entrytime="00:00:24.50" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="10305" heatid="10730" lane="5" entrytime="00:02:18.00" />
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="10306" heatid="10751" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="10307" heatid="10817" lane="9" entrytime="00:01:20.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="10308" heatid="10838" lane="4" entrytime="00:00:25.00" />
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="10309" heatid="10904" lane="5" entrytime="00:02:20.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="10310" heatid="10925" lane="6" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Hubert" gender="M" lastname="Markowski" nation="POL" athleteid="9682">
              <RESULTS>
                <RESULT eventid="1190" points="350" swimtime="00:02:41.64" resultid="9922" heatid="10727" lane="1" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:14.68" />
                    <SPLIT distance="150" swimtime="00:02:03.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="340" swimtime="00:00:34.41" resultid="9923" heatid="10748" lane="8" entrytime="00:00:34.50" />
                <RESULT eventid="1452" points="333" swimtime="00:01:14.75" resultid="9924" heatid="10847" lane="4" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="323" swimtime="00:05:55.19" resultid="9925" heatid="10879" lane="4" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:14.89" />
                    <SPLIT distance="150" swimtime="00:02:02.96" />
                    <SPLIT distance="200" swimtime="00:02:49.54" />
                    <SPLIT distance="250" swimtime="00:03:40.27" />
                    <SPLIT distance="300" swimtime="00:04:32.19" />
                    <SPLIT distance="350" swimtime="00:05:15.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Piotr" gender="M" lastname="Biankowski" nation="POL" athleteid="7227">
              <RESULTS>
                <RESULT eventid="1128" points="254" swimtime="00:22:54.04" resultid="10277" heatid="10677" lane="2" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                    <SPLIT distance="100" swimtime="00:01:25.72" />
                    <SPLIT distance="150" swimtime="00:02:11.95" />
                    <SPLIT distance="200" swimtime="00:02:57.37" />
                    <SPLIT distance="250" swimtime="00:03:42.81" />
                    <SPLIT distance="300" swimtime="00:04:29.06" />
                    <SPLIT distance="350" swimtime="00:05:14.54" />
                    <SPLIT distance="400" swimtime="00:06:00.26" />
                    <SPLIT distance="450" swimtime="00:06:45.72" />
                    <SPLIT distance="500" swimtime="00:07:31.77" />
                    <SPLIT distance="550" swimtime="00:08:18.01" />
                    <SPLIT distance="600" swimtime="00:09:04.54" />
                    <SPLIT distance="650" swimtime="00:09:50.77" />
                    <SPLIT distance="700" swimtime="00:10:37.44" />
                    <SPLIT distance="750" swimtime="00:11:23.55" />
                    <SPLIT distance="800" swimtime="00:12:10.00" />
                    <SPLIT distance="850" swimtime="00:12:56.20" />
                    <SPLIT distance="900" swimtime="00:13:42.83" />
                    <SPLIT distance="950" swimtime="00:14:28.81" />
                    <SPLIT distance="1000" swimtime="00:15:15.44" />
                    <SPLIT distance="1050" swimtime="00:16:01.62" />
                    <SPLIT distance="1100" swimtime="00:16:48.07" />
                    <SPLIT distance="1150" swimtime="00:17:34.08" />
                    <SPLIT distance="1200" swimtime="00:18:20.61" />
                    <SPLIT distance="1250" swimtime="00:19:06.45" />
                    <SPLIT distance="1300" swimtime="00:19:52.56" />
                    <SPLIT distance="1350" swimtime="00:20:38.93" />
                    <SPLIT distance="1400" swimtime="00:21:25.27" />
                    <SPLIT distance="1450" swimtime="00:22:10.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="259" swimtime="00:02:58.63" resultid="10278" heatid="10721" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:26.63" />
                    <SPLIT distance="150" swimtime="00:02:20.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="216" swimtime="00:03:05.57" resultid="10279" heatid="10794" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:25.05" />
                    <SPLIT distance="150" swimtime="00:02:13.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" status="DNS" swimtime="00:00:00.00" resultid="10280" heatid="10878" lane="0" entrytime="00:07:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Piotr" gender="M" lastname="Koliński" nation="POL" athleteid="10653">
              <RESULTS>
                <RESULT eventid="1160" points="320" swimtime="00:00:30.54" resultid="10654" heatid="10698" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1302" points="299" swimtime="00:01:10.14" resultid="10655" heatid="10779" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="291" swimtime="00:00:33.82" resultid="10656" heatid="10830" lane="7" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Zbigniew" gender="M" lastname="Paluszak" nation="POL" athleteid="7277">
              <RESULTS>
                <RESULT eventid="1160" points="85" swimtime="00:00:47.48" resultid="9808" heatid="10691" lane="0" entrytime="00:00:47.85" />
                <RESULT eventid="1302" points="83" swimtime="00:01:47.31" resultid="9809" heatid="10773" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="104" swimtime="00:02:01.47" resultid="9810" heatid="10809" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="149" swimtime="00:00:49.73" resultid="9811" heatid="10913" lane="4" entrytime="00:00:52.35" />
                <RESULT eventid="1695" points="88" swimtime="00:08:14.01" resultid="9812" heatid="10935" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.18" />
                    <SPLIT distance="100" swimtime="00:01:49.29" />
                    <SPLIT distance="150" swimtime="00:02:53.34" />
                    <SPLIT distance="200" swimtime="00:03:57.80" />
                    <SPLIT distance="250" swimtime="00:05:01.17" />
                    <SPLIT distance="300" swimtime="00:06:06.48" />
                    <SPLIT distance="350" swimtime="00:07:10.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Janusz" gender="M" lastname="Płonka" nation="POL" athleteid="9835">
              <RESULTS>
                <RESULT eventid="1190" points="56" swimtime="00:04:56.43" resultid="9836" heatid="10719" lane="4" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.55" />
                    <SPLIT distance="100" swimtime="00:02:26.10" />
                    <SPLIT distance="150" swimtime="00:03:59.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="88" swimtime="00:00:53.98" resultid="9837" heatid="10741" lane="5" entrytime="00:00:56.00" />
                <RESULT eventid="1332" points="41" swimtime="00:05:23.19" resultid="9838" heatid="10791" lane="5" entrytime="00:05:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.06" />
                    <SPLIT distance="100" swimtime="00:02:31.94" />
                    <SPLIT distance="150" swimtime="00:04:02.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="96" swimtime="00:00:48.95" resultid="9839" heatid="10826" lane="6" entrytime="00:00:52.00" />
                <RESULT eventid="1546" points="52" swimtime="00:10:50.98" resultid="9840" heatid="10876" lane="2" entrytime="00:10:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.88" />
                    <SPLIT distance="100" swimtime="00:02:26.93" />
                    <SPLIT distance="150" swimtime="00:04:03.58" />
                    <SPLIT distance="200" swimtime="00:05:28.65" />
                    <SPLIT distance="250" swimtime="00:07:00.57" />
                    <SPLIT distance="300" swimtime="00:08:31.36" />
                    <SPLIT distance="350" swimtime="00:09:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="47" swimtime="00:02:17.11" resultid="9841" heatid="10885" lane="6" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="49" swimtime="00:10:00.71" resultid="9842" heatid="10936" lane="1" entrytime="00:09:22.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:03:42.52" />
                    <SPLIT distance="200" swimtime="00:05:05.34" />
                    <SPLIT distance="250" swimtime="00:06:23.43" />
                    <SPLIT distance="350" swimtime="00:07:15.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Petr" gender="M" lastname="HORVÁT" nation="POL" athleteid="10643">
              <RESULTS>
                <RESULT eventid="1160" points="484" swimtime="00:00:26.63" resultid="10644" heatid="10708" lane="2" entrytime="00:00:26.60" />
                <RESULT eventid="1190" points="481" swimtime="00:02:25.46" resultid="10645" heatid="10730" lane="7" entrytime="00:02:23.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:08.95" />
                    <SPLIT distance="150" swimtime="00:01:52.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="445" swimtime="00:00:31.48" resultid="10646" heatid="10750" lane="5" entrytime="00:00:30.87" />
                <RESULT eventid="1332" points="403" swimtime="00:02:30.87" resultid="10647" heatid="10796" lane="7" entrytime="00:02:29.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                    <SPLIT distance="150" swimtime="00:01:51.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="485" swimtime="00:01:05.95" resultid="10648" heatid="10849" lane="4" entrytime="00:01:06.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="468" swimtime="00:05:13.97" resultid="10649" heatid="10881" lane="1" entrytime="00:05:12.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:13.85" />
                    <SPLIT distance="150" swimtime="00:01:52.32" />
                    <SPLIT distance="200" swimtime="00:02:32.26" />
                    <SPLIT distance="250" swimtime="00:03:17.25" />
                    <SPLIT distance="300" swimtime="00:04:03.69" />
                    <SPLIT distance="350" swimtime="00:04:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="447" swimtime="00:02:26.28" resultid="10650" heatid="10904" lane="3" entrytime="00:02:25.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                    <SPLIT distance="100" swimtime="00:01:11.56" />
                    <SPLIT distance="150" swimtime="00:01:49.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="475" swimtime="00:04:41.87" resultid="10651" heatid="10945" lane="8" entrytime="00:04:40.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                    <SPLIT distance="100" swimtime="00:01:05.97" />
                    <SPLIT distance="150" swimtime="00:01:42.45" />
                    <SPLIT distance="200" swimtime="00:02:18.57" />
                    <SPLIT distance="250" swimtime="00:02:55.04" />
                    <SPLIT distance="300" swimtime="00:03:31.36" />
                    <SPLIT distance="350" swimtime="00:04:07.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Krzysztof" gender="M" lastname="Drózd" nation="POL" athleteid="9760">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="9909" heatid="10705" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="1242" points="353" swimtime="00:00:34.00" resultid="9910" heatid="10747" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="373" swimtime="00:01:05.12" resultid="9911" heatid="10781" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="290" swimtime="00:01:18.26" resultid="9912" heatid="10847" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="291" swimtime="00:02:33.82" resultid="9913" heatid="10861" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:01:53.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="9914" heatid="10902" lane="4" entrytime="00:02:45.00" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="9915" heatid="10938" lane="4" entrytime="00:06:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Bolesław" gender="M" lastname="Czyż" nation="POL" athleteid="6208" />
            <ATHLETE birthdate="1987-01-01" firstname="Dorota" gender="F" lastname="Szczypiór" nation="POL" athleteid="7297">
              <RESULTS>
                <RESULT eventid="1144" points="364" swimtime="00:00:33.23" resultid="10318" heatid="10681" lane="8" />
                <RESULT eventid="1175" points="229" swimtime="00:03:25.88" resultid="10319" heatid="10712" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                    <SPLIT distance="100" swimtime="00:01:38.69" />
                    <SPLIT distance="150" swimtime="00:02:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="297" swimtime="00:01:17.96" resultid="10320" heatid="10765" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Krzysztof" gender="M" lastname="Kępa" nation="POL" athleteid="6221">
              <RESULTS>
                <RESULT eventid="1160" points="247" swimtime="00:00:33.32" resultid="10568" heatid="10696" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="231" swimtime="00:01:16.45" resultid="10569" heatid="10775" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="10570" heatid="10858" lane="5" entrytime="00:03:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="6231">
              <RESULTS>
                <RESULT eventid="1160" points="388" swimtime="00:00:28.66" resultid="10576" heatid="10704" lane="9" entrytime="00:00:28.75" />
                <RESULT eventid="1190" points="337" swimtime="00:02:43.79" resultid="10577" heatid="10726" lane="6" entrytime="00:02:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:16.91" />
                    <SPLIT distance="150" swimtime="00:02:07.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="393" swimtime="00:01:04.03" resultid="10578" heatid="10782" lane="2" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="383" swimtime="00:00:30.86" resultid="10579" heatid="10833" lane="2" entrytime="00:00:30.85" />
                <RESULT eventid="1452" points="286" swimtime="00:01:18.63" resultid="10580" heatid="10848" lane="1" entrytime="00:01:15.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="332" swimtime="00:01:11.88" resultid="10581" heatid="10889" lane="2" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="330" swimtime="00:00:38.22" resultid="10582" heatid="10921" lane="0" entrytime="00:00:37.75" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Leandro" gender="M" lastname="Pascua" nation="POL" athleteid="7195">
              <RESULTS>
                <RESULT eventid="1332" status="DNS" swimtime="00:00:00.00" resultid="10260" heatid="10794" lane="8" entrytime="00:03:05.00" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="10261" heatid="10942" lane="3" entrytime="00:05:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Yauheni" gender="M" lastname="Puzan" nation="POL" athleteid="7283">
              <RESULTS>
                <RESULT eventid="1160" points="559" swimtime="00:00:25.37" resultid="10311" heatid="10710" lane="5" entrytime="00:00:25.00" />
                <RESULT eventid="1242" points="603" swimtime="00:00:28.45" resultid="10312" heatid="10751" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1302" points="619" swimtime="00:00:55.04" resultid="10313" heatid="10788" lane="6" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="698" swimtime="00:00:25.28" resultid="10314" heatid="10838" lane="3" entrytime="00:00:25.50" />
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="10315" heatid="10863" lane="1" entrytime="00:02:20.00" />
                <RESULT eventid="1578" points="649" swimtime="00:00:57.53" resultid="10316" heatid="10892" lane="4" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="439" swimtime="00:00:34.75" resultid="10317" heatid="10923" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Piotr" gender="M" lastname="Krzekotowski" nation="POL" athleteid="7236">
              <RESULTS>
                <RESULT eventid="1160" points="160" swimtime="00:00:38.47" resultid="10281" heatid="10693" lane="9" entrytime="00:00:39.01" />
                <RESULT eventid="1190" points="113" swimtime="00:03:55.65" resultid="10282" heatid="10719" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.83" />
                    <SPLIT distance="100" swimtime="00:02:03.31" />
                    <SPLIT distance="150" swimtime="00:03:07.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="129" swimtime="00:04:11.22" resultid="10283" heatid="10758" lane="0" entrytime="00:04:15.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.39" />
                    <SPLIT distance="100" swimtime="00:02:00.02" />
                    <SPLIT distance="150" swimtime="00:03:05.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="139" swimtime="00:01:30.46" resultid="10284" heatid="10774" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="108" swimtime="00:01:59.80" resultid="10285" heatid="10810" lane="3" entrytime="00:01:51.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="115" swimtime="00:03:29.60" resultid="10286" heatid="10857" lane="3" entrytime="00:03:29.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.62" />
                    <SPLIT distance="100" swimtime="00:01:38.36" />
                    <SPLIT distance="150" swimtime="00:02:34.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Konrad" gender="M" lastname="Szydło" nation="POL" athleteid="9747">
              <RESULTS>
                <RESULT eventid="1128" points="269" swimtime="00:22:28.35" resultid="10946" heatid="10677" lane="5" late="yes" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:17.50" />
                    <SPLIT distance="150" swimtime="00:01:59.94" />
                    <SPLIT distance="200" swimtime="00:02:44.57" />
                    <SPLIT distance="250" swimtime="00:03:28.28" />
                    <SPLIT distance="300" swimtime="00:04:13.43" />
                    <SPLIT distance="350" swimtime="00:04:57.94" />
                    <SPLIT distance="400" swimtime="00:05:42.89" />
                    <SPLIT distance="450" swimtime="00:06:26.70" />
                    <SPLIT distance="500" swimtime="00:07:12.05" />
                    <SPLIT distance="550" swimtime="00:07:55.48" />
                    <SPLIT distance="600" swimtime="00:08:40.28" />
                    <SPLIT distance="650" swimtime="00:09:24.38" />
                    <SPLIT distance="700" swimtime="00:10:09.82" />
                    <SPLIT distance="750" swimtime="00:10:55.08" />
                    <SPLIT distance="800" swimtime="00:11:41.08" />
                    <SPLIT distance="850" swimtime="00:12:26.61" />
                    <SPLIT distance="900" swimtime="00:13:13.58" />
                    <SPLIT distance="950" swimtime="00:14:00.19" />
                    <SPLIT distance="1000" swimtime="00:14:47.11" />
                    <SPLIT distance="1050" swimtime="00:15:33.57" />
                    <SPLIT distance="1100" swimtime="00:16:20.37" />
                    <SPLIT distance="1150" swimtime="00:17:07.19" />
                    <SPLIT distance="1200" swimtime="00:17:54.08" />
                    <SPLIT distance="1250" swimtime="00:18:41.22" />
                    <SPLIT distance="1300" swimtime="00:19:28.83" />
                    <SPLIT distance="1350" swimtime="00:20:14.40" />
                    <SPLIT distance="1400" swimtime="00:21:00.30" />
                    <SPLIT distance="1450" swimtime="00:21:45.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="340" swimtime="00:00:29.95" resultid="10947" heatid="10701" lane="4" late="yes" entrytime="00:00:29.59" />
                <RESULT eventid="1242" points="277" swimtime="00:00:36.87" resultid="10948" heatid="10747" lane="7" entrytime="00:00:35.30" />
                <RESULT eventid="1302" points="340" swimtime="00:01:07.18" resultid="10949" heatid="10780" lane="3" entrytime="00:01:06.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="278" swimtime="00:01:19.41" resultid="10950" heatid="10847" lane="2" entrytime="00:01:19.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="298" swimtime="00:02:32.61" resultid="10951" heatid="10861" lane="3" entrytime="00:02:28.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="150" swimtime="00:01:54.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="271" swimtime="00:02:52.88" resultid="10952" heatid="10902" lane="1" entrytime="00:02:56.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                    <SPLIT distance="150" swimtime="00:02:09.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="10953" heatid="10941" lane="4" entrytime="00:05:20.36" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="7205">
              <RESULTS>
                <RESULT eventid="1128" points="208" swimtime="00:24:29.02" resultid="10265" heatid="10676" lane="9" entrytime="00:25:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                    <SPLIT distance="100" swimtime="00:01:30.23" />
                    <SPLIT distance="150" swimtime="00:02:18.58" />
                    <SPLIT distance="200" swimtime="00:03:09.11" />
                    <SPLIT distance="250" swimtime="00:03:57.84" />
                    <SPLIT distance="300" swimtime="00:04:47.18" />
                    <SPLIT distance="350" swimtime="00:05:36.70" />
                    <SPLIT distance="400" swimtime="00:06:25.54" />
                    <SPLIT distance="450" swimtime="00:07:14.51" />
                    <SPLIT distance="500" swimtime="00:08:03.85" />
                    <SPLIT distance="550" swimtime="00:08:53.22" />
                    <SPLIT distance="600" swimtime="00:09:43.80" />
                    <SPLIT distance="650" swimtime="00:10:33.42" />
                    <SPLIT distance="700" swimtime="00:11:23.76" />
                    <SPLIT distance="750" swimtime="00:12:14.03" />
                    <SPLIT distance="800" swimtime="00:13:03.36" />
                    <SPLIT distance="850" swimtime="00:13:52.41" />
                    <SPLIT distance="900" swimtime="00:14:42.83" />
                    <SPLIT distance="950" swimtime="00:15:33.24" />
                    <SPLIT distance="1000" swimtime="00:16:22.08" />
                    <SPLIT distance="1050" swimtime="00:17:11.01" />
                    <SPLIT distance="1100" swimtime="00:18:01.50" />
                    <SPLIT distance="1150" swimtime="00:18:51.14" />
                    <SPLIT distance="1200" swimtime="00:19:39.94" />
                    <SPLIT distance="1250" swimtime="00:20:24.43" />
                    <SPLIT distance="1300" swimtime="00:21:18.81" />
                    <SPLIT distance="1350" swimtime="00:22:08.02" />
                    <SPLIT distance="1400" swimtime="00:22:56.41" />
                    <SPLIT distance="1450" swimtime="00:23:45.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="275" swimtime="00:00:32.13" resultid="10266" heatid="10697" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1302" points="267" swimtime="00:01:12.76" resultid="10267" heatid="10778" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="10268" heatid="10828" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1482" points="203" swimtime="00:02:53.30" resultid="10269" heatid="10859" lane="6" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                    <SPLIT distance="150" swimtime="00:02:09.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="10270" heatid="10915" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1695" points="209" swimtime="00:06:10.68" resultid="10271" heatid="10939" lane="0" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:27.13" />
                    <SPLIT distance="150" swimtime="00:02:15.79" />
                    <SPLIT distance="200" swimtime="00:03:04.45" />
                    <SPLIT distance="250" swimtime="00:03:53.13" />
                    <SPLIT distance="300" swimtime="00:04:41.82" />
                    <SPLIT distance="350" swimtime="00:05:28.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Andrii" gender="M" lastname="Moraru" nation="POL" athleteid="7271">
              <RESULTS>
                <RESULT eventid="1160" points="227" swimtime="00:00:34.26" resultid="9818" heatid="10694" lane="2" entrytime="00:00:35.92" />
                <RESULT eventid="1242" points="125" swimtime="00:00:48.01" resultid="9819" heatid="10742" lane="6" entrytime="00:00:51.10" />
                <RESULT eventid="1392" points="193" swimtime="00:01:38.77" resultid="9820" heatid="10812" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="119" swimtime="00:00:45.58" resultid="9821" heatid="10827" lane="8" entrytime="00:00:46.08" />
                <RESULT eventid="1638" points="210" swimtime="00:00:44.38" resultid="9822" heatid="10916" lane="0" entrytime="00:00:43.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Bernard" gender="M" lastname="Filek" nation="POL" athleteid="9506">
              <RESULTS>
                <RESULT eventid="1160" points="521" swimtime="00:00:25.97" resultid="10954" heatid="10710" lane="0" late="yes" entrytime="00:00:25.50" />
                <RESULT eventid="1242" points="448" swimtime="00:00:31.41" resultid="10955" heatid="10751" lane="6" late="yes" entrytime="00:00:30.00" />
                <RESULT eventid="1302" points="549" swimtime="00:00:57.26" resultid="10956" heatid="10788" lane="7" late="yes" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="549" swimtime="00:00:27.39" resultid="10957" heatid="10837" lane="4" late="yes" entrytime="00:00:27.00" />
                <RESULT eventid="1452" points="386" swimtime="00:01:11.18" resultid="10958" heatid="10843" lane="7" late="yes" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Paweł" gender="M" lastname="Borkowski" nation="POL" athleteid="7201">
              <RESULTS>
                <RESULT eventid="1160" points="420" swimtime="00:00:27.90" resultid="10262" heatid="10702" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1302" points="465" swimtime="00:01:00.55" resultid="10263" heatid="10782" lane="8" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="10264" heatid="10861" lane="2" entrytime="00:02:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Paweł" gender="M" lastname="Marudzinski" nation="POL" athleteid="6216">
              <RESULTS>
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="10564" heatid="10671" lane="5" entrytime="00:11:29.91" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="10565" heatid="10761" lane="6" entrytime="00:03:05.90" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="10566" heatid="10815" lane="3" entrytime="00:01:24.05" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="10567" heatid="10921" lane="9" entrytime="00:00:37.84" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Luca" gender="M" lastname="Manfredi" nation="POL" athleteid="7249">
              <RESULTS>
                <RESULT eventid="1160" points="562" swimtime="00:00:25.33" resultid="10292" heatid="10711" lane="9" entrytime="00:00:24.90" />
                <RESULT eventid="1302" points="548" swimtime="00:00:57.30" resultid="10293" heatid="10787" lane="5" entrytime="00:00:55.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Joanna" gender="F" lastname="Matysiak" nation="POL" athleteid="9215">
              <RESULTS>
                <RESULT eventid="1144" points="364" swimtime="00:00:33.22" resultid="11060" heatid="10681" lane="9" late="yes" />
                <RESULT eventid="1226" status="DNS" swimtime="00:00:00.00" resultid="11061" heatid="10734" lane="9" late="yes" />
                <RESULT eventid="1376" points="237" swimtime="00:01:43.88" resultid="11062" heatid="10803" lane="8" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="228" swimtime="00:01:35.01" resultid="11063" heatid="10839" lane="9" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Adrianna" gender="F" lastname="Buraczynska" nation="POL" athleteid="6202">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="10553" heatid="10667" lane="1" entrytime="00:13:00.00" />
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="10554" heatid="10717" lane="8" entrytime="00:02:55.00" />
                <RESULT eventid="1226" points="510" swimtime="00:00:33.86" resultid="10555" heatid="10738" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1437" points="474" swimtime="00:01:14.51" resultid="10556" heatid="10842" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="410" swimtime="00:02:46.91" resultid="10557" heatid="10897" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="100" swimtime="00:01:19.79" />
                    <SPLIT distance="150" swimtime="00:02:03.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Aleksandra" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="10297">
              <RESULTS>
                <RESULT eventid="1144" points="521" swimtime="00:00:29.48" resultid="10298" heatid="10688" lane="0" entrytime="00:00:29.50" />
                <RESULT eventid="1226" points="516" swimtime="00:00:33.72" resultid="10299" heatid="10739" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1287" status="DNS" swimtime="00:00:00.00" resultid="10300" heatid="10770" lane="6" entrytime="00:01:09.50" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="10301" heatid="10842" lane="7" entrytime="00:01:14.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="Michał" gender="M" lastname="Mandes" nation="POL" athleteid="10641">
              <RESULTS>
                <RESULT eventid="1422" points="402" swimtime="00:00:30.39" resultid="10642" heatid="10834" lane="5" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-04-09" firstname="Anna" gender="F" lastname="Błazucka" nation="POL" athleteid="7539">
              <RESULTS>
                <RESULT eventid="1144" points="76" swimtime="00:00:55.81" resultid="10605" heatid="10681" lane="6" entrytime="00:00:56.40" entrycourse="SCM" />
                <RESULT eventid="1226" points="45" swimtime="00:01:15.69" resultid="10606" heatid="10734" lane="1" />
                <RESULT eventid="1257" points="62" swimtime="00:05:50.28" resultid="10607" heatid="10753" lane="9" entrytime="00:05:27.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.78" />
                    <SPLIT distance="100" swimtime="00:02:48.68" />
                    <SPLIT distance="150" swimtime="00:04:21.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="52" swimtime="00:02:52.21" resultid="10608" heatid="10803" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="58" swimtime="00:01:16.08" resultid="10609" heatid="10905" lane="4" entrytime="00:01:12.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-01-01" firstname="Andrzej" gender="M" lastname="Deptuła" nation="POL" athleteid="11054">
              <RESULTS>
                <RESULT eventid="1160" points="15" swimtime="00:01:24.05" resultid="11055" heatid="10691" lane="9" late="yes" />
                <RESULT eventid="1302" points="6" swimtime="00:04:11.25" resultid="11056" heatid="10772" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:54.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="11057" heatid="10825" lane="6" late="yes" />
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="11058" heatid="10856" lane="0" late="yes" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="11059" heatid="10885" lane="9" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Kazimierz" gender="M" lastname="Sinicki" nation="POL" athleteid="7232">
              <RESULTS>
                <RESULT eventid="1160" points="315" swimtime="00:00:30.72" resultid="9926" heatid="10699" lane="1" entrytime="00:00:31.15" />
                <RESULT eventid="1302" points="299" swimtime="00:01:10.10" resultid="9927" heatid="10778" lane="5" entrytime="00:01:10.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="230" swimtime="00:02:46.33" resultid="9928" heatid="10860" lane="7" entrytime="00:02:45.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                    <SPLIT distance="150" swimtime="00:02:02.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Mateusz" gender="M" lastname="Dymiter" nation="POL" athleteid="9794">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="9795" heatid="10697" lane="9" entrytime="00:00:33.00" />
                <RESULT comment="G 8 - Ukończenie wyścigu nie w położeniu na plecach" eventid="1190" status="DSQ" swimtime="00:02:38.66" resultid="9796" heatid="10724" lane="4" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:15.43" />
                    <SPLIT distance="150" swimtime="00:02:01.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="311" swimtime="00:00:35.46" resultid="9797" heatid="10746" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1302" points="373" swimtime="00:01:05.14" resultid="9798" heatid="10777" lane="8" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="314" swimtime="00:01:23.98" resultid="9799" heatid="10812" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="290" swimtime="00:01:18.31" resultid="9800" heatid="10846" lane="5" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="367" swimtime="00:01:09.58" resultid="9801" heatid="10887" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="311" swimtime="00:00:38.96" resultid="9802" heatid="10919" lane="9" entrytime="00:00:39.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Maciej" gender="M" lastname="Lubas" nation="POL" athleteid="7243">
              <RESULTS>
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="10287" heatid="10669" lane="1" entrytime="00:23:30.00" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="10288" heatid="10726" lane="9" entrytime="00:02:47.00" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="10289" heatid="10763" lane="0" entrytime="00:02:50.00" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="10290" heatid="10817" lane="8" entrytime="00:01:18.50" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="10291" heatid="10924" lane="9" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Tomasz" gender="M" lastname="Ciesielski" nation="POL" athleteid="9773">
              <RESULTS>
                <RESULT eventid="1160" points="418" swimtime="00:00:27.96" resultid="9828" heatid="10705" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1190" points="289" swimtime="00:02:52.30" resultid="9829" heatid="10729" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:14.68" />
                    <SPLIT distance="150" swimtime="00:02:06.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="9830" heatid="10750" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="9831" heatid="10834" lane="9" entrytime="00:00:30.50" />
                <RESULT eventid="1452" status="DNS" swimtime="00:00:00.00" resultid="9832" heatid="10848" lane="5" entrytime="00:01:12.00" />
                <RESULT eventid="1608" points="262" swimtime="00:02:54.79" resultid="9833" heatid="10904" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:01:19.56" />
                    <SPLIT distance="150" swimtime="00:02:07.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="417" swimtime="00:00:35.36" resultid="9834" heatid="10922" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-11" firstname="Paweł" gender="M" lastname="Adamowicz" nation="POL" athleteid="7101">
              <RESULTS>
                <RESULT eventid="1160" points="139" swimtime="00:00:40.35" resultid="9787" heatid="10692" lane="9" entrytime="00:00:42.16" entrycourse="LCM" />
                <RESULT eventid="1392" points="183" swimtime="00:01:40.60" resultid="9788" heatid="10811" lane="7" entrytime="00:01:45.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="215" swimtime="00:00:44.08" resultid="9789" heatid="10915" lane="4" entrytime="00:00:44.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Petr" gender="M" lastname="Horvát" nation="POL" athleteid="10251">
              <RESULTS>
                <RESULT eventid="1160" points="291" swimtime="00:00:31.53" resultid="10252" heatid="10700" lane="3" entrytime="00:00:30.11" />
                <RESULT eventid="1190" points="244" swimtime="00:03:02.28" resultid="10253" heatid="10722" lane="4" entrytime="00:03:08.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:30.51" />
                    <SPLIT distance="150" swimtime="00:02:22.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="200" swimtime="00:00:41.05" resultid="10254" heatid="10745" lane="6" entrytime="00:00:39.32" />
                <RESULT eventid="1272" points="310" swimtime="00:03:07.63" resultid="10255" heatid="10761" lane="3" entrytime="00:03:05.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="100" swimtime="00:01:31.22" />
                    <SPLIT distance="150" swimtime="00:02:19.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="295" swimtime="00:01:25.82" resultid="10256" heatid="10815" lane="9" entrytime="00:01:26.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="253" swimtime="00:02:41.16" resultid="10257" heatid="10860" lane="2" entrytime="00:02:44.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                    <SPLIT distance="100" swimtime="00:01:17.25" />
                    <SPLIT distance="150" swimtime="00:02:00.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="186" swimtime="00:01:27.15" resultid="10258" heatid="10887" lane="9" entrytime="00:01:30.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="318" swimtime="00:00:38.69" resultid="10259" heatid="10920" lane="4" entrytime="00:00:37.87" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEKRA" nation="POL" region="MAŁ" clubid="3166" name="Niezrzeszony Kraków">
          <CONTACT email="piotr_urbanczyk@onet.pl" name="URBAŃCZYK PIOTR" phone="608172201" />
          <ATHLETES>
            <ATHLETE birthdate="1984-03-16" firstname="Piotr" gender="M" lastname="Urbańczyk" nation="POL" athleteid="6600">
              <RESULTS>
                <RESULT eventid="1242" points="509" swimtime="00:00:30.09" resultid="6601" heatid="10751" lane="1" entrytime="00:00:28.99" />
                <RESULT eventid="1452" points="517" swimtime="00:01:04.59" resultid="6602" heatid="10850" lane="4" entrytime="00:01:02.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="471" swimtime="00:02:23.81" resultid="6603" heatid="10904" lane="4" entrytime="00:02:19.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                    <SPLIT distance="150" swimtime="00:01:47.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIERAD" nation="POL" region="14" clubid="6175" name="Niezrzeszony Radom">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1953-01-01" firstname="Wlodzimierz" gender="M" lastname="Zieleziński" nation="POL" athleteid="6239">
              <RESULTS>
                <RESULT eventid="1160" points="222" swimtime="00:00:34.52" resultid="7525" heatid="10695" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1242" points="184" swimtime="00:00:42.26" resultid="7526" heatid="10744" lane="3" entrytime="00:00:41.50" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="7527" heatid="10777" lane="0" entrytime="00:01:18.00" />
                <RESULT eventid="1452" points="144" swimtime="00:01:38.71" resultid="7528" heatid="10845" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="7529" heatid="10858" lane="2" entrytime="00:03:03.00" />
                <RESULT eventid="1608" points="138" swimtime="00:03:36.36" resultid="7530" heatid="10900" lane="6" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.47" />
                    <SPLIT distance="100" swimtime="00:01:45.86" />
                    <SPLIT distance="150" swimtime="00:02:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="7531" heatid="10938" lane="2" entrytime="00:06:25.00" />
                <RESULT eventid="1128" status="DNS" swimtime="00:00:00.00" resultid="9516" heatid="10675" lane="6" entrytime="00:26:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEZR1" nation="POL" region="14" clubid="9929" name="Niezrzeszony1">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Konrad" gender="M" lastname="Jajecznik" nation="POL" athleteid="10658">
              <RESULTS>
                <RESULT eventid="1160" points="141" swimtime="00:00:40.15" resultid="10659" heatid="10692" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1302" points="142" swimtime="00:01:29.77" resultid="10660" heatid="10774" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="139" swimtime="00:00:43.20" resultid="10661" heatid="10827" lane="9" entrytime="00:00:47.00" />
                <RESULT eventid="1482" points="137" swimtime="00:03:17.84" resultid="10662" heatid="10857" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:01:33.97" />
                    <SPLIT distance="150" swimtime="00:02:26.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="232" swimtime="00:00:42.94" resultid="10663" heatid="10918" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1695" points="145" swimtime="00:06:58.32" resultid="10664" heatid="10936" lane="6" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                    <SPLIT distance="100" swimtime="00:01:34.63" />
                    <SPLIT distance="150" swimtime="00:02:25.70" />
                    <SPLIT distance="200" swimtime="00:03:21.39" />
                    <SPLIT distance="250" swimtime="00:04:16.42" />
                    <SPLIT distance="300" swimtime="00:05:12.32" />
                    <SPLIT distance="350" swimtime="00:06:07.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Marcin" gender="M" lastname="Warda" nation="POL" athleteid="9987">
              <RESULTS>
                <RESULT eventid="1160" points="277" swimtime="00:00:32.05" resultid="10039" heatid="10698" lane="2" entrytime="00:00:31.75" />
                <RESULT eventid="1638" points="259" swimtime="00:00:41.42" resultid="10040" heatid="10917" lane="3" entrytime="00:00:40.48" />
                <RESULT eventid="1695" points="186" swimtime="00:06:25.20" resultid="10041" heatid="10938" lane="3" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:14.05" />
                    <SPLIT distance="200" swimtime="00:03:03.73" />
                    <SPLIT distance="250" swimtime="00:03:54.85" />
                    <SPLIT distance="300" swimtime="00:04:46.37" />
                    <SPLIT distance="350" swimtime="00:05:38.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEZR2" nation="POL" region="14" clubid="10052" name="Niezrzeszony2">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1977-01-01" firstname="Marek" gender="M" lastname="Gizicki" nation="POL" athleteid="10109">
              <RESULTS>
                <RESULT eventid="1128" points="232" swimtime="00:23:35.86" resultid="10110" heatid="10677" lane="9" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                    <SPLIT distance="100" swimtime="00:01:23.17" />
                    <SPLIT distance="150" swimtime="00:02:08.45" />
                    <SPLIT distance="200" swimtime="00:02:54.29" />
                    <SPLIT distance="250" swimtime="00:03:41.10" />
                    <SPLIT distance="300" swimtime="00:04:28.28" />
                    <SPLIT distance="350" swimtime="00:05:16.28" />
                    <SPLIT distance="400" swimtime="00:06:03.98" />
                    <SPLIT distance="450" swimtime="00:06:51.87" />
                    <SPLIT distance="500" swimtime="00:07:39.82" />
                    <SPLIT distance="550" swimtime="00:08:28.11" />
                    <SPLIT distance="600" swimtime="00:09:16.21" />
                    <SPLIT distance="650" swimtime="00:10:04.80" />
                    <SPLIT distance="700" swimtime="00:10:52.54" />
                    <SPLIT distance="750" swimtime="00:11:40.83" />
                    <SPLIT distance="800" swimtime="00:12:28.81" />
                    <SPLIT distance="850" swimtime="00:13:17.37" />
                    <SPLIT distance="900" swimtime="00:14:05.25" />
                    <SPLIT distance="950" swimtime="00:14:54.19" />
                    <SPLIT distance="1000" swimtime="00:15:41.93" />
                    <SPLIT distance="1050" swimtime="00:16:30.04" />
                    <SPLIT distance="1100" swimtime="00:17:18.01" />
                    <SPLIT distance="1150" swimtime="00:18:07.52" />
                    <SPLIT distance="1200" swimtime="00:18:55.78" />
                    <SPLIT distance="1250" swimtime="00:19:44.40" />
                    <SPLIT distance="1300" swimtime="00:20:32.24" />
                    <SPLIT distance="1350" swimtime="00:21:20.45" />
                    <SPLIT distance="1400" swimtime="00:22:07.10" />
                    <SPLIT distance="1450" swimtime="00:22:40.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Alan" gender="M" lastname="Bistron" nation="POL" athleteid="10090">
              <RESULTS>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="10091" heatid="10898" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Magdaena" gender="F" lastname="Jezierska" nation="POL" athleteid="10085">
              <RESULTS>
                <RESULT eventid="1175" points="283" swimtime="00:03:12.02" resultid="10086" heatid="10715" lane="0" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="150" swimtime="00:02:21.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="401" swimtime="00:00:36.67" resultid="10087" heatid="10738" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1407" points="281" swimtime="00:00:37.28" resultid="10088" heatid="10823" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1437" points="366" swimtime="00:01:21.20" resultid="10089" heatid="10841" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Jolanta" gender="F" lastname="Zawadzka" nation="POL" athleteid="10092">
              <RESULTS>
                <RESULT eventid="1175" points="208" swimtime="00:03:32.86" resultid="10093" heatid="10714" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                    <SPLIT distance="100" swimtime="00:01:41.43" />
                    <SPLIT distance="150" swimtime="00:02:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="261" swimtime="00:01:40.57" resultid="10094" heatid="10805" lane="6" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="213" swimtime="00:00:40.86" resultid="10095" heatid="10821" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1623" points="270" swimtime="00:00:45.59" resultid="10096" heatid="10908" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Dorota" gender="F" lastname="Batóg" nation="POL" athleteid="10102">
              <RESULTS>
                <RESULT eventid="1144" points="329" swimtime="00:00:34.34" resultid="10103" heatid="10685" lane="1" entrytime="00:00:34.35" />
                <RESULT eventid="1226" points="250" swimtime="00:00:42.92" resultid="10104" heatid="10737" lane="7" entrytime="00:00:41.73" />
                <RESULT eventid="1287" points="278" swimtime="00:01:19.76" resultid="10105" heatid="10768" lane="2" entrytime="00:01:19.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="267" swimtime="00:01:39.93" resultid="10106" heatid="10805" lane="3" entrytime="00:01:41.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="205" swimtime="00:00:41.39" resultid="10107" heatid="10822" lane="0" entrytime="00:00:39.35" />
                <RESULT eventid="1623" points="294" swimtime="00:00:44.32" resultid="10108" heatid="10908" lane="5" entrytime="00:00:44.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Wiesław" gender="M" lastname="Bar" nation="POL" athleteid="10078">
              <RESULTS>
                <RESULT eventid="1128" points="316" swimtime="00:21:18.29" resultid="10079" heatid="10678" lane="4" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="150" swimtime="00:01:54.20" />
                    <SPLIT distance="200" swimtime="00:02:35.82" />
                    <SPLIT distance="250" swimtime="00:03:17.34" />
                    <SPLIT distance="300" swimtime="00:03:59.53" />
                    <SPLIT distance="350" swimtime="00:04:42.02" />
                    <SPLIT distance="400" swimtime="00:05:24.49" />
                    <SPLIT distance="450" swimtime="00:06:07.47" />
                    <SPLIT distance="500" swimtime="00:06:50.49" />
                    <SPLIT distance="550" swimtime="00:07:33.84" />
                    <SPLIT distance="600" swimtime="00:08:17.44" />
                    <SPLIT distance="650" swimtime="00:09:01.33" />
                    <SPLIT distance="700" swimtime="00:09:44.60" />
                    <SPLIT distance="750" swimtime="00:10:28.10" />
                    <SPLIT distance="800" swimtime="00:11:11.67" />
                    <SPLIT distance="850" swimtime="00:11:55.73" />
                    <SPLIT distance="900" swimtime="00:12:39.82" />
                    <SPLIT distance="950" swimtime="00:13:23.80" />
                    <SPLIT distance="1000" swimtime="00:14:07.53" />
                    <SPLIT distance="1050" swimtime="00:14:51.33" />
                    <SPLIT distance="1100" swimtime="00:15:34.88" />
                    <SPLIT distance="1150" swimtime="00:16:18.83" />
                    <SPLIT distance="1200" swimtime="00:17:02.59" />
                    <SPLIT distance="1250" swimtime="00:17:46.33" />
                    <SPLIT distance="1300" swimtime="00:18:29.88" />
                    <SPLIT distance="1350" swimtime="00:19:13.51" />
                    <SPLIT distance="1400" swimtime="00:19:56.38" />
                    <SPLIT distance="1450" swimtime="00:20:39.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="390" swimtime="00:00:28.61" resultid="10080" heatid="10705" lane="9" entrytime="00:00:28.00" />
                <RESULT eventid="1190" points="333" swimtime="00:02:44.44" resultid="10081" heatid="10726" lane="2" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:02:07.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="343" swimtime="00:00:34.33" resultid="10082" heatid="10748" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1302" points="396" swimtime="00:01:03.85" resultid="10083" heatid="10783" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="10084" heatid="10863" lane="4" entrytime="00:02:17.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NOSTA" nation="UKR" clubid="5008" name="NoStars">
          <CONTACT email="nostarsswimming@gmail.com" internet="www.nostarsclub.ru" name="Krot Stanislav" phone="+38 050 4651785" zip="14000" />
          <ATHLETES>
            <ATHLETE birthdate="1962-08-09" firstname="Igor" gender="M" lastname="Medvediev" nation="UKR" athleteid="5009">
              <RESULTS>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="7545" heatid="10729" lane="9" entrytime="00:02:33.00" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="7546" heatid="10763" lane="2" entrytime="00:02:47.00" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="7547" heatid="10818" lane="3" entrytime="00:01:14.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="7548" heatid="10925" lane="0" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AQODE" nation="UKR" clubid="5014" name="Odessa Aqua Masters">
          <CONTACT email="imedvedev99@rambler.ru" name="Medvediev Igor" phone="+38 050 7866547" />
          <ATHLETES>
            <ATHLETE birthdate="1952-12-12" firstname="Dymytrii" gender="M" lastname="Malinovskyi" nation="UKR" athleteid="5015">
              <RESULTS>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="7556" heatid="10758" lane="5" entrytime="00:03:45.00" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="7557" heatid="10813" lane="0" entrytime="00:01:35.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="7558" heatid="10886" lane="2" entrytime="00:01:42.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="7559" heatid="10917" lane="1" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MATAR" nation="POL" region="SLA" clubid="5267" name="Park Wodny Tarnowskie Góry Masters Team" shortname="Park Wodny Tarnowskie Góry Mas">
          <CONTACT city="Tarnowskie Góry" email="swimman@o2.pl" name="Pąchalski Tomasz" phone="600-365-944" state="SLA" street="Obwodnica 8" zip="42-600" />
          <ATHLETES>
            <ATHLETE birthdate="1975-08-09" firstname="Sonia" gender="F" lastname="Borkowska" nation="POL" athleteid="5273">
              <RESULTS>
                <RESULT eventid="1144" points="367" swimtime="00:00:33.14" resultid="8291" heatid="10686" lane="7" entrytime="00:00:33.05" />
                <RESULT eventid="1287" points="327" swimtime="00:01:15.56" resultid="8292" heatid="10769" lane="7" entrytime="00:01:15.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="237" swimtime="00:01:43.85" resultid="8293" heatid="10806" lane="5" entrytime="00:01:35.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="265" swimtime="00:02:55.79" resultid="8294" heatid="10854" lane="6" entrytime="00:02:45.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                    <SPLIT distance="100" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:02:09.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PLKAI" nation="LTU" clubid="2913" name="Plaukiam Kaisaidorys">
          <CONTACT city="Vilnius" email="alex@gedwood.eu" name="Aleksandras" phone="+370 65609220" street="Fiziku 14-59" zip="VNO" />
          <ATHLETES>
            <ATHLETE birthdate="1971-04-22" firstname="Aleksandras" gender="M" lastname="Zamorskis" nation="LTU" athleteid="2914">
              <RESULTS>
                <RESULT eventid="1190" points="509" swimtime="00:02:22.72" resultid="7781" heatid="10730" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                    <SPLIT distance="100" swimtime="00:01:06.96" />
                    <SPLIT distance="150" swimtime="00:01:48.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="521" swimtime="00:00:58.29" resultid="7782" heatid="10787" lane="9" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="497" swimtime="00:00:28.31" resultid="7783" heatid="10836" lane="7" entrytime="00:00:28.50" />
                <RESULT eventid="1482" points="464" swimtime="00:02:11.74" resultid="7784" heatid="10865" lane="3" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:01:04.89" />
                    <SPLIT distance="150" swimtime="00:01:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="439" swimtime="00:01:05.53" resultid="7785" heatid="10891" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="551" swimtime="00:00:32.22" resultid="7786" heatid="10925" lane="5" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-19" firstname="Eimantas" gender="M" lastname="Frankonis" nation="LTU" athleteid="2921">
              <RESULTS>
                <RESULT eventid="1272" points="308" swimtime="00:03:08.05" resultid="7787" heatid="10762" lane="7" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                    <SPLIT distance="100" swimtime="00:01:27.87" />
                    <SPLIT distance="150" swimtime="00:02:17.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="336" swimtime="00:01:22.13" resultid="7788" heatid="10816" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="356" swimtime="00:00:37.26" resultid="7789" heatid="10922" lane="7" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-07-20" firstname="Raimondas" gender="M" lastname="Gincas" nation="LTU" athleteid="2930">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="7794" heatid="10708" lane="5" entrytime="00:00:26.50" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="7795" heatid="10786" lane="7" entrytime="00:00:59.00" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="7796" heatid="10817" lane="6" entrytime="00:01:17.00" />
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="7797" heatid="10864" lane="1" entrytime="00:02:15.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="7798" heatid="10922" lane="5" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-17" firstname="Mantas" gender="M" lastname="Petrulis" nation="LTU" athleteid="2925">
              <RESULTS>
                <RESULT eventid="1160" points="451" swimtime="00:00:27.25" resultid="7790" heatid="10707" lane="2" entrytime="00:00:27.00" />
                <RESULT eventid="1392" points="412" swimtime="00:01:16.74" resultid="7791" heatid="10818" lane="9" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="462" swimtime="00:00:29.01" resultid="7792" heatid="10836" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1638" points="497" swimtime="00:00:33.34" resultid="7793" heatid="10925" lane="8" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1518" status="DNS" swimtime="00:00:00.00" resultid="7799" heatid="10871" lane="4" entrytime="00:01:53.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2914" number="1" />
                    <RELAYPOSITION athleteid="2925" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2921" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2930" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1368" status="DNS" swimtime="00:00:00.00" resultid="7800" heatid="10802" lane="8" entrytime="00:02:02.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2914" number="1" />
                    <RELAYPOSITION athleteid="2921" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2925" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2930" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SLPL" nation="CZE" clubid="3390" name="Plavecký klub Slávia VŠ Plzeň">
          <CONTACT city="Plzeň" email="srailova@bazenslovany.cz" internet="www.bazenslovany.cz/plavecky-klub" name="Radka Bažilová" state="CZE" street="náměstí Generála Píky 42" zip="32600" />
          <ATHLETES>
            <ATHLETE birthdate="1946-05-17" firstname="Petr" gender="M" lastname="Buble" nation="CZE" athleteid="5202">
              <RESULTS>
                <RESULT eventid="1272" points="240" swimtime="00:03:24.24" resultid="7830" heatid="10760" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.70" />
                    <SPLIT distance="100" swimtime="00:01:37.96" />
                    <SPLIT distance="150" swimtime="00:02:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="230" swimtime="00:01:33.22" resultid="7831" heatid="10813" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="193" swimtime="00:03:13.39" resultid="7832" heatid="10901" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                    <SPLIT distance="100" swimtime="00:01:35.32" />
                    <SPLIT distance="150" swimtime="00:02:24.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-10-18" firstname="Kamila" gender="F" lastname="Častoral" nation="CZE" athleteid="5206">
              <RESULTS>
                <RESULT eventid="1257" points="144" swimtime="00:04:24.97" resultid="7833" heatid="10754" lane="0" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.53" />
                    <SPLIT distance="100" swimtime="00:02:10.48" />
                    <SPLIT distance="150" swimtime="00:03:18.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="147" swimtime="00:02:01.81" resultid="7834" heatid="10804" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="167" swimtime="00:00:53.53" resultid="7835" heatid="10907" lane="2" entrytime="00:00:50.00" />
                <RESULT comment="M 7 - Nieprzenoszenie ramion do przodu nad lustrem wody" eventid="1525" status="DSQ" swimtime="00:09:38.99" resultid="9654" heatid="10873" lane="6" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.62" />
                    <SPLIT distance="100" swimtime="00:02:29.77" />
                    <SPLIT distance="150" swimtime="00:03:51.44" />
                    <SPLIT distance="200" swimtime="00:05:06.42" />
                    <SPLIT distance="250" swimtime="00:06:15.05" />
                    <SPLIT distance="300" swimtime="00:07:22.36" />
                    <SPLIT distance="350" swimtime="00:08:31.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="85" swimtime="00:04:41.09" resultid="9655" heatid="10894" lane="7" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.80" />
                    <SPLIT distance="100" swimtime="00:02:22.51" />
                    <SPLIT distance="150" swimtime="00:03:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="90" swimtime="00:04:40.63" resultid="9823" heatid="10713" lane="8" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.97" />
                    <SPLIT distance="100" swimtime="00:02:22.75" />
                    <SPLIT distance="150" swimtime="00:03:33.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-06-07" firstname="Daniel" gender="M" lastname="Štěpán" nation="CZE" athleteid="5198">
              <RESULTS>
                <RESULT eventid="1302" points="296" swimtime="00:01:10.33" resultid="7827" heatid="10776" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="233" swimtime="00:02:45.69" resultid="7828" heatid="10858" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:17.28" />
                    <SPLIT distance="150" swimtime="00:02:02.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="216" swimtime="00:06:06.75" resultid="7829" heatid="10939" lane="8" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:23.24" />
                    <SPLIT distance="150" swimtime="00:02:09.87" />
                    <SPLIT distance="200" swimtime="00:02:57.96" />
                    <SPLIT distance="250" swimtime="00:03:46.45" />
                    <SPLIT distance="300" swimtime="00:04:35.02" />
                    <SPLIT distance="350" swimtime="00:05:23.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TEOGR" nation="POL" region="14" clubid="6185" name="Polish Ogrodnik Team">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Bogusław" gender="M" lastname="Ogrodnik" nation="POL" athleteid="6248">
              <RESULTS>
                <RESULT eventid="1128" points="152" swimtime="00:27:11.23" resultid="7533" heatid="10676" lane="2" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:01:33.07" />
                    <SPLIT distance="150" swimtime="00:02:23.91" />
                    <SPLIT distance="200" swimtime="00:03:17.14" />
                    <SPLIT distance="250" swimtime="00:04:11.27" />
                    <SPLIT distance="300" swimtime="00:05:04.85" />
                    <SPLIT distance="350" swimtime="00:05:59.14" />
                    <SPLIT distance="400" swimtime="00:06:53.59" />
                    <SPLIT distance="450" swimtime="00:07:48.96" />
                    <SPLIT distance="500" swimtime="00:08:44.39" />
                    <SPLIT distance="550" swimtime="00:09:39.25" />
                    <SPLIT distance="600" swimtime="00:10:35.22" />
                    <SPLIT distance="650" swimtime="00:11:31.09" />
                    <SPLIT distance="700" swimtime="00:12:26.43" />
                    <SPLIT distance="750" swimtime="00:13:21.21" />
                    <SPLIT distance="800" swimtime="00:14:16.99" />
                    <SPLIT distance="850" swimtime="00:15:12.44" />
                    <SPLIT distance="900" swimtime="00:16:09.13" />
                    <SPLIT distance="950" swimtime="00:17:05.45" />
                    <SPLIT distance="1000" swimtime="00:18:00.31" />
                    <SPLIT distance="1050" swimtime="00:18:57.51" />
                    <SPLIT distance="1100" swimtime="00:19:53.00" />
                    <SPLIT distance="1150" swimtime="00:20:48.80" />
                    <SPLIT distance="1200" swimtime="00:21:43.89" />
                    <SPLIT distance="1250" swimtime="00:22:39.59" />
                    <SPLIT distance="1300" swimtime="00:23:36.20" />
                    <SPLIT distance="1350" swimtime="00:24:31.71" />
                    <SPLIT distance="1400" swimtime="00:25:25.96" />
                    <SPLIT distance="1450" swimtime="00:26:20.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="183" swimtime="00:00:36.82" resultid="7534" heatid="10696" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1302" points="208" swimtime="00:01:19.16" resultid="7535" heatid="10777" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="158" swimtime="00:01:45.57" resultid="7536" heatid="10811" lane="5" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="163" swimtime="00:03:06.55" resultid="7537" heatid="10859" lane="0" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:25.89" />
                    <SPLIT distance="150" swimtime="00:02:17.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PRKAL" nation="RUS" clubid="5825" name="Pregel Kaliningrad">
          <CONTACT name="s" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Vadim" gender="M" lastname="Ezhkov" nation="RUS" athleteid="5913">
              <RESULTS>
                <RESULT eventid="1128" points="279" swimtime="00:22:12.83" resultid="7402" heatid="10678" lane="2" entrytime="00:21:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="150" swimtime="00:02:02.18" />
                    <SPLIT distance="200" swimtime="00:02:45.82" />
                    <SPLIT distance="250" swimtime="00:03:29.45" />
                    <SPLIT distance="300" swimtime="00:04:13.36" />
                    <SPLIT distance="350" swimtime="00:04:57.39" />
                    <SPLIT distance="400" swimtime="00:05:41.71" />
                    <SPLIT distance="450" swimtime="00:06:26.18" />
                    <SPLIT distance="500" swimtime="00:07:11.00" />
                    <SPLIT distance="550" swimtime="00:07:54.70" />
                    <SPLIT distance="600" swimtime="00:08:39.41" />
                    <SPLIT distance="650" swimtime="00:09:23.89" />
                    <SPLIT distance="700" swimtime="00:10:09.14" />
                    <SPLIT distance="750" swimtime="00:10:53.74" />
                    <SPLIT distance="800" swimtime="00:11:38.92" />
                    <SPLIT distance="850" swimtime="00:12:23.71" />
                    <SPLIT distance="900" swimtime="00:13:09.38" />
                    <SPLIT distance="950" swimtime="00:13:54.07" />
                    <SPLIT distance="1000" swimtime="00:14:39.76" />
                    <SPLIT distance="1050" swimtime="00:15:24.96" />
                    <SPLIT distance="1100" swimtime="00:16:11.32" />
                    <SPLIT distance="1150" swimtime="00:16:56.59" />
                    <SPLIT distance="1200" swimtime="00:17:42.89" />
                    <SPLIT distance="1250" swimtime="00:18:27.86" />
                    <SPLIT distance="1300" swimtime="00:19:13.82" />
                    <SPLIT distance="1350" swimtime="00:19:59.35" />
                    <SPLIT distance="1400" swimtime="00:20:45.79" />
                    <SPLIT distance="1450" swimtime="00:21:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="291" swimtime="00:00:31.53" resultid="7403" heatid="10700" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1190" points="270" swimtime="00:02:56.23" resultid="7404" heatid="10724" lane="6" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:27.56" />
                    <SPLIT distance="150" swimtime="00:02:16.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="297" swimtime="00:01:25.54" resultid="7405" heatid="10815" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="211" swimtime="00:01:27.05" resultid="7406" heatid="10846" lane="8" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="358" swimtime="00:00:37.19" resultid="7407" heatid="10921" lane="8" entrytime="00:00:37.50" />
                <RESULT eventid="1695" points="294" swimtime="00:05:30.94" resultid="7408" heatid="10941" lane="2" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:18.71" />
                    <SPLIT distance="150" swimtime="00:02:01.31" />
                    <SPLIT distance="200" swimtime="00:02:44.61" />
                    <SPLIT distance="250" swimtime="00:03:26.59" />
                    <SPLIT distance="300" swimtime="00:04:10.02" />
                    <SPLIT distance="350" swimtime="00:04:51.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Elena" gender="F" lastname="Koliadyna" nation="RUS" athleteid="5831">
              <RESULTS>
                <RESULT eventid="1144" points="285" swimtime="00:00:36.02" resultid="7334" heatid="10684" lane="4" entrytime="00:00:35.50" />
                <RESULT eventid="1257" points="256" swimtime="00:03:38.93" resultid="7335" heatid="10754" lane="5" entrytime="00:03:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.20" />
                    <SPLIT distance="100" swimtime="00:01:44.33" />
                    <SPLIT distance="150" swimtime="00:02:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="247" swimtime="00:01:42.44" resultid="7336" heatid="10806" lane="8" entrytime="00:01:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.79" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O 9 - Przepłynięcie przez zawodnika na inny tor podczas wyścigu" eventid="1437" status="DSQ" swimtime="00:01:50.83" resultid="7337" heatid="10840" lane="7" entrytime="00:01:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="302" swimtime="00:00:43.92" resultid="7338" heatid="10908" lane="3" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Viacheslav" gender="M" lastname="Tikhonov" nation="RUS" athleteid="5879">
              <RESULTS>
                <RESULT eventid="1160" points="194" swimtime="00:00:36.06" resultid="7374" heatid="10694" lane="6" entrytime="00:00:35.50" />
                <RESULT eventid="1242" points="140" swimtime="00:00:46.25" resultid="7375" heatid="10743" lane="7" entrytime="00:00:46.50" />
                <RESULT eventid="1422" points="124" swimtime="00:00:44.98" resultid="7376" heatid="10827" lane="7" entrytime="00:00:45.50" />
                <RESULT eventid="1638" points="158" swimtime="00:00:48.84" resultid="7377" heatid="10915" lane="0" entrytime="00:00:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Oksana" gender="F" lastname="Bronitskaya" nation="RUS" athleteid="5855">
              <RESULTS>
                <RESULT eventid="1175" points="499" swimtime="00:02:38.92" resultid="7354" heatid="10718" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="150" swimtime="00:02:01.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="456" swimtime="00:00:35.14" resultid="7355" heatid="10739" lane="1" entrytime="00:00:34.50" />
                <RESULT eventid="1257" points="452" swimtime="00:03:01.21" resultid="7356" heatid="10756" lane="6" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:27.51" />
                    <SPLIT distance="150" swimtime="00:02:14.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="447" swimtime="00:00:31.93" resultid="7357" heatid="10824" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="1525" points="447" swimtime="00:05:48.32" resultid="7358" heatid="10875" lane="3" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:06.57" />
                    <SPLIT distance="200" swimtime="00:02:54.01" />
                    <SPLIT distance="250" swimtime="00:03:41.86" />
                    <SPLIT distance="300" swimtime="00:04:32.22" />
                    <SPLIT distance="350" swimtime="00:05:10.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="425" swimtime="00:02:44.91" resultid="7359" heatid="10897" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:01:20.73" />
                    <SPLIT distance="150" swimtime="00:02:02.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="447" swimtime="00:05:09.09" resultid="7360" heatid="10934" lane="2" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:01:54.56" />
                    <SPLIT distance="200" swimtime="00:02:34.21" />
                    <SPLIT distance="250" swimtime="00:03:13.99" />
                    <SPLIT distance="300" swimtime="00:03:53.64" />
                    <SPLIT distance="350" swimtime="00:04:31.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-01-01" firstname="Luiza" gender="F" lastname="Shcherbich" nation="RUS" athleteid="5826">
              <RESULTS>
                <RESULT eventid="1144" points="49" swimtime="00:01:04.83" resultid="7330" heatid="10681" lane="7" entrytime="00:01:05.00" />
                <RESULT eventid="1257" points="64" swimtime="00:05:46.93" resultid="7331" heatid="10752" lane="4" entrytime="00:05:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.52" />
                    <SPLIT distance="100" swimtime="00:02:57.81" />
                    <SPLIT distance="150" swimtime="00:04:27.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="51" swimtime="00:02:53.34" resultid="7332" heatid="10803" lane="6" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="61" swimtime="00:01:14.86" resultid="7333" heatid="10905" lane="5" entrytime="00:01:13.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-01" firstname="Aleksandr" gender="M" lastname="Tervinskii" nation="RUS" athleteid="5898">
              <RESULTS>
                <RESULT eventid="1160" points="217" swimtime="00:00:34.76" resultid="7390" heatid="10695" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1242" points="171" swimtime="00:00:43.27" resultid="7391" heatid="10744" lane="0" entrytime="00:00:42.80" />
                <RESULT eventid="1392" points="167" swimtime="00:01:43.67" resultid="7392" heatid="10811" lane="3" entrytime="00:01:42.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="239" swimtime="00:00:42.56" resultid="7393" heatid="10916" lane="2" entrytime="00:00:42.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Regina" gender="F" lastname="Sych" nation="RUS" athleteid="5873">
              <RESULTS>
                <RESULT eventid="1144" points="657" swimtime="00:00:27.29" resultid="7369" heatid="10688" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="1287" points="655" swimtime="00:00:59.92" resultid="7370" heatid="10771" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="563" swimtime="00:00:29.57" resultid="7371" heatid="10824" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="1467" points="576" swimtime="00:02:15.72" resultid="7372" heatid="10855" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:05.84" />
                    <SPLIT distance="150" swimtime="00:01:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" status="DNS" swimtime="00:00:00.00" resultid="7373" heatid="10934" lane="3" entrytime="00:04:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Aleksandr" gender="M" lastname="Smirnov" nation="RUS" athleteid="5921">
              <RESULTS>
                <RESULT eventid="1128" points="390" swimtime="00:19:51.92" resultid="7409" heatid="10679" lane="2" entrytime="00:19:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:52.52" />
                    <SPLIT distance="200" swimtime="00:02:32.12" />
                    <SPLIT distance="250" swimtime="00:03:11.06" />
                    <SPLIT distance="300" swimtime="00:03:50.44" />
                    <SPLIT distance="350" swimtime="00:04:29.45" />
                    <SPLIT distance="400" swimtime="00:05:08.98" />
                    <SPLIT distance="450" swimtime="00:05:47.81" />
                    <SPLIT distance="500" swimtime="00:06:27.25" />
                    <SPLIT distance="550" swimtime="00:07:06.64" />
                    <SPLIT distance="600" swimtime="00:07:46.41" />
                    <SPLIT distance="650" swimtime="00:08:26.63" />
                    <SPLIT distance="700" swimtime="00:09:06.76" />
                    <SPLIT distance="750" swimtime="00:09:46.65" />
                    <SPLIT distance="800" swimtime="00:10:27.26" />
                    <SPLIT distance="850" swimtime="00:11:07.03" />
                    <SPLIT distance="900" swimtime="00:11:47.74" />
                    <SPLIT distance="950" swimtime="00:12:27.61" />
                    <SPLIT distance="1000" swimtime="00:13:08.46" />
                    <SPLIT distance="1050" swimtime="00:13:45.39" />
                    <SPLIT distance="1100" swimtime="00:14:29.70" />
                    <SPLIT distance="1150" swimtime="00:15:10.69" />
                    <SPLIT distance="1200" swimtime="00:15:51.76" />
                    <SPLIT distance="1250" swimtime="00:16:16.74" />
                    <SPLIT distance="1350" swimtime="00:16:32.41" />
                    <SPLIT distance="1400" swimtime="00:17:13.18" />
                    <SPLIT distance="1450" swimtime="00:17:53.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="7410" heatid="10703" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="7411" heatid="10782" lane="5" entrytime="00:01:03.50" />
                <RESULT eventid="1482" points="380" swimtime="00:02:20.72" resultid="7412" heatid="10863" lane="6" entrytime="00:02:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:46.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="399" swimtime="00:04:58.89" resultid="7413" heatid="10943" lane="6" entrytime="00:05:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:11.01" />
                    <SPLIT distance="150" swimtime="00:01:49.24" />
                    <SPLIT distance="200" swimtime="00:02:27.75" />
                    <SPLIT distance="250" swimtime="00:03:06.27" />
                    <SPLIT distance="300" swimtime="00:03:44.52" />
                    <SPLIT distance="350" swimtime="00:04:22.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Yuri" gender="M" lastname="Yakovenko" nation="RUS" athleteid="5884">
              <RESULTS>
                <RESULT eventid="1160" points="168" swimtime="00:00:37.89" resultid="7378" heatid="10693" lane="5" entrytime="00:00:37.50" />
                <RESULT eventid="1272" points="147" swimtime="00:04:00.57" resultid="7379" heatid="10758" lane="2" entrytime="00:03:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.67" />
                    <SPLIT distance="100" swimtime="00:01:57.52" />
                    <SPLIT distance="150" swimtime="00:03:00.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="155" swimtime="00:01:46.31" resultid="7380" heatid="10811" lane="0" entrytime="00:01:47.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="193" swimtime="00:00:45.64" resultid="7381" heatid="10915" lane="7" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Eduard" gender="M" lastname="Bersenev" nation="RUS" athleteid="5889">
              <RESULTS>
                <RESULT eventid="1160" points="243" swimtime="00:00:33.50" resultid="7382" heatid="10700" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1190" points="208" swimtime="00:03:12.22" resultid="7383" heatid="10723" lane="4" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="100" swimtime="00:01:34.43" />
                    <SPLIT distance="150" swimtime="00:02:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="201" swimtime="00:00:41.02" resultid="7384" heatid="10745" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1302" points="268" swimtime="00:01:12.67" resultid="7385" heatid="10778" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="260" swimtime="00:00:35.12" resultid="7386" heatid="10830" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1482" points="252" swimtime="00:02:41.41" resultid="7387" heatid="10860" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                    <SPLIT distance="100" swimtime="00:01:18.43" />
                    <SPLIT distance="150" swimtime="00:02:00.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="215" swimtime="00:00:44.05" resultid="7388" heatid="10916" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1695" points="247" swimtime="00:05:50.36" resultid="7389" heatid="10940" lane="7" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                    <SPLIT distance="100" swimtime="00:01:21.78" />
                    <SPLIT distance="150" swimtime="00:02:06.53" />
                    <SPLIT distance="200" swimtime="00:02:51.36" />
                    <SPLIT distance="250" swimtime="00:03:37.01" />
                    <SPLIT distance="300" swimtime="00:04:21.93" />
                    <SPLIT distance="350" swimtime="00:05:07.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Irina" gender="F" lastname="Titova" nation="RUS" athleteid="5850">
              <RESULTS>
                <RESULT eventid="1144" points="300" swimtime="00:00:35.43" resultid="7350" heatid="10685" lane="9" entrytime="00:00:35.50" />
                <RESULT eventid="1287" points="320" swimtime="00:01:16.04" resultid="7351" heatid="10769" lane="8" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="314" swimtime="00:02:46.11" resultid="7352" heatid="10854" lane="7" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:19.76" />
                    <SPLIT distance="150" swimtime="00:02:03.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="304" swimtime="00:05:51.48" resultid="7353" heatid="10933" lane="5" entrytime="00:05:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:23.16" />
                    <SPLIT distance="150" swimtime="00:02:08.30" />
                    <SPLIT distance="200" swimtime="00:02:53.68" />
                    <SPLIT distance="250" swimtime="00:03:38.96" />
                    <SPLIT distance="300" swimtime="00:04:24.34" />
                    <SPLIT distance="350" swimtime="00:05:09.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Sergei" gender="M" lastname="Karakchiev" nation="RUS" athleteid="5927">
              <RESULTS>
                <RESULT eventid="1160" points="398" swimtime="00:00:28.42" resultid="7414" heatid="10706" lane="0" entrytime="00:00:27.50" />
                <RESULT eventid="1242" points="397" swimtime="00:00:32.69" resultid="7415" heatid="10748" lane="3" entrytime="00:00:33.50" />
                <RESULT eventid="1452" points="379" swimtime="00:01:11.61" resultid="7416" heatid="10848" lane="3" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="337" swimtime="00:02:40.78" resultid="7417" heatid="10903" lane="1" entrytime="00:02:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:16.93" />
                    <SPLIT distance="150" swimtime="00:01:57.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Liudmila" gender="F" lastname="Kokhan" nation="RUS" athleteid="5868">
              <RESULTS>
                <RESULT eventid="1144" points="365" swimtime="00:00:33.20" resultid="7365" heatid="10685" lane="8" entrytime="00:00:34.80" />
                <RESULT eventid="1287" points="299" swimtime="00:01:17.80" resultid="7366" heatid="10768" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="263" swimtime="00:01:40.41" resultid="7367" heatid="10805" lane="8" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="268" swimtime="00:00:45.68" resultid="7368" heatid="10907" lane="3" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Sergei" gender="M" lastname="Mikhaylov" nation="RUS" athleteid="5903">
              <RESULTS>
                <RESULT eventid="1128" points="172" swimtime="00:26:05.44" resultid="7394" heatid="10675" lane="8" entrytime="00:30:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.62" />
                    <SPLIT distance="100" swimtime="00:01:36.61" />
                    <SPLIT distance="150" swimtime="00:02:28.64" />
                    <SPLIT distance="200" swimtime="00:03:20.43" />
                    <SPLIT distance="250" swimtime="00:04:12.91" />
                    <SPLIT distance="300" swimtime="00:05:04.77" />
                    <SPLIT distance="350" swimtime="00:05:57.45" />
                    <SPLIT distance="400" swimtime="00:06:48.78" />
                    <SPLIT distance="450" swimtime="00:07:40.11" />
                    <SPLIT distance="500" swimtime="00:08:31.69" />
                    <SPLIT distance="550" swimtime="00:09:24.18" />
                    <SPLIT distance="600" swimtime="00:10:16.34" />
                    <SPLIT distance="650" swimtime="00:11:09.09" />
                    <SPLIT distance="700" swimtime="00:12:02.01" />
                    <SPLIT distance="750" swimtime="00:12:54.70" />
                    <SPLIT distance="800" swimtime="00:13:47.59" />
                    <SPLIT distance="850" swimtime="00:14:40.39" />
                    <SPLIT distance="900" swimtime="00:15:33.91" />
                    <SPLIT distance="950" swimtime="00:16:26.99" />
                    <SPLIT distance="1000" swimtime="00:17:20.32" />
                    <SPLIT distance="1050" swimtime="00:18:12.84" />
                    <SPLIT distance="1100" swimtime="00:19:06.29" />
                    <SPLIT distance="1150" swimtime="00:19:59.26" />
                    <SPLIT distance="1200" swimtime="00:20:53.20" />
                    <SPLIT distance="1250" swimtime="00:21:46.72" />
                    <SPLIT distance="1300" swimtime="00:22:39.83" />
                    <SPLIT distance="1350" swimtime="00:23:32.46" />
                    <SPLIT distance="1400" swimtime="00:24:25.71" />
                    <SPLIT distance="1450" swimtime="00:25:16.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Natalia" gender="F" lastname="Aleshchenko" nation="RUS" athleteid="5837">
              <RESULTS>
                <RESULT eventid="1113" points="251" swimtime="00:24:26.40" resultid="7339" heatid="10674" lane="2" entrytime="00:24:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                    <SPLIT distance="100" swimtime="00:01:28.93" />
                    <SPLIT distance="150" swimtime="00:02:16.91" />
                    <SPLIT distance="200" swimtime="00:03:04.57" />
                    <SPLIT distance="250" swimtime="00:03:52.09" />
                    <SPLIT distance="300" swimtime="00:04:39.66" />
                    <SPLIT distance="350" swimtime="00:05:27.81" />
                    <SPLIT distance="400" swimtime="00:06:15.43" />
                    <SPLIT distance="450" swimtime="00:07:03.58" />
                    <SPLIT distance="500" swimtime="00:07:50.85" />
                    <SPLIT distance="550" swimtime="00:08:39.15" />
                    <SPLIT distance="600" swimtime="00:09:27.11" />
                    <SPLIT distance="650" swimtime="00:10:16.16" />
                    <SPLIT distance="700" swimtime="00:11:04.62" />
                    <SPLIT distance="750" swimtime="00:11:54.37" />
                    <SPLIT distance="800" swimtime="00:12:43.23" />
                    <SPLIT distance="850" swimtime="00:13:33.03" />
                    <SPLIT distance="900" swimtime="00:14:22.88" />
                    <SPLIT distance="950" swimtime="00:15:13.80" />
                    <SPLIT distance="1000" swimtime="00:16:03.49" />
                    <SPLIT distance="1050" swimtime="00:16:54.49" />
                    <SPLIT distance="1100" swimtime="00:17:44.55" />
                    <SPLIT distance="1150" swimtime="00:18:35.57" />
                    <SPLIT distance="1200" swimtime="00:19:26.03" />
                    <SPLIT distance="1250" swimtime="00:20:17.75" />
                    <SPLIT distance="1300" swimtime="00:21:08.25" />
                    <SPLIT distance="1350" swimtime="00:21:59.51" />
                    <SPLIT distance="1400" swimtime="00:22:50.37" />
                    <SPLIT distance="1450" swimtime="00:23:41.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="278" swimtime="00:03:13.18" resultid="7340" heatid="10715" lane="9" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                    <SPLIT distance="100" swimtime="00:01:35.25" />
                    <SPLIT distance="150" swimtime="00:02:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="215" swimtime="00:00:45.14" resultid="7341" heatid="10736" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1287" points="272" swimtime="00:01:20.29" resultid="7342" heatid="10768" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="245" swimtime="00:00:39.04" resultid="7343" heatid="10822" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="1467" points="267" swimtime="00:02:55.39" resultid="7344" heatid="10854" lane="8" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                    <SPLIT distance="100" swimtime="00:01:26.16" />
                    <SPLIT distance="150" swimtime="00:02:12.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="194" swimtime="00:03:34.07" resultid="7345" heatid="10895" lane="0" entrytime="00:03:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.09" />
                    <SPLIT distance="100" swimtime="00:01:46.01" />
                    <SPLIT distance="150" swimtime="00:02:41.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="267" swimtime="00:06:07.14" resultid="7346" heatid="10933" lane="1" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                    <SPLIT distance="100" swimtime="00:01:28.15" />
                    <SPLIT distance="150" swimtime="00:02:16.06" />
                    <SPLIT distance="200" swimtime="00:03:03.98" />
                    <SPLIT distance="250" swimtime="00:03:51.60" />
                    <SPLIT distance="300" swimtime="00:04:39.20" />
                    <SPLIT distance="350" swimtime="00:05:25.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Grigorii" gender="M" lastname="Lopin" nation="RUS" athleteid="5905">
              <RESULTS>
                <RESULT eventid="1098" points="237" swimtime="00:12:09.58" resultid="7395" heatid="10671" lane="8" entrytime="00:11:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                    <SPLIT distance="100" swimtime="00:01:21.22" />
                    <SPLIT distance="150" swimtime="00:02:07.17" />
                    <SPLIT distance="200" swimtime="00:02:54.07" />
                    <SPLIT distance="250" swimtime="00:03:41.38" />
                    <SPLIT distance="300" swimtime="00:04:28.03" />
                    <SPLIT distance="350" swimtime="00:05:14.88" />
                    <SPLIT distance="400" swimtime="00:06:02.53" />
                    <SPLIT distance="450" swimtime="00:06:48.23" />
                    <SPLIT distance="500" swimtime="00:07:34.05" />
                    <SPLIT distance="550" swimtime="00:08:20.83" />
                    <SPLIT distance="600" swimtime="00:09:07.97" />
                    <SPLIT distance="650" swimtime="00:09:54.99" />
                    <SPLIT distance="700" swimtime="00:10:41.32" />
                    <SPLIT distance="750" swimtime="00:11:27.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="299" swimtime="00:00:31.26" resultid="7396" heatid="10699" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1272" points="267" swimtime="00:03:17.18" resultid="7397" heatid="10760" lane="3" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                    <SPLIT distance="100" swimtime="00:01:36.55" />
                    <SPLIT distance="150" swimtime="00:02:27.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="279" swimtime="00:01:27.42" resultid="7398" heatid="10814" lane="0" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="225" swimtime="00:06:40.37" resultid="7399" heatid="10878" lane="7" entrytime="00:06:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.39" />
                    <SPLIT distance="100" swimtime="00:01:38.75" />
                    <SPLIT distance="150" swimtime="00:02:33.42" />
                    <SPLIT distance="200" swimtime="00:03:28.30" />
                    <SPLIT distance="250" swimtime="00:04:20.25" />
                    <SPLIT distance="300" swimtime="00:05:13.49" />
                    <SPLIT distance="350" swimtime="00:05:56.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="298" swimtime="00:00:39.52" resultid="7400" heatid="10919" lane="0" entrytime="00:00:39.50" />
                <RESULT eventid="1695" points="234" swimtime="00:05:56.79" resultid="7401" heatid="10940" lane="4" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.52" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:08.68" />
                    <SPLIT distance="200" swimtime="00:02:55.76" />
                    <SPLIT distance="250" swimtime="00:03:42.33" />
                    <SPLIT distance="300" swimtime="00:04:28.75" />
                    <SPLIT distance="350" swimtime="00:05:15.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Liudmila" gender="F" lastname="Skopina" nation="RUS" athleteid="5846">
              <RESULTS>
                <RESULT eventid="1257" points="189" swimtime="00:04:02.32" resultid="7347" heatid="10753" lane="4" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.27" />
                    <SPLIT distance="100" swimtime="00:01:57.42" />
                    <SPLIT distance="150" swimtime="00:03:00.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="195" swimtime="00:01:50.94" resultid="7348" heatid="10804" lane="5" entrytime="00:01:51.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="208" swimtime="00:00:49.73" resultid="7349" heatid="10907" lane="1" entrytime="00:00:51.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="201" swimtime="00:02:39.38" resultid="7431" heatid="10800" lane="2" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.31" />
                    <SPLIT distance="100" swimtime="00:01:27.30" />
                    <SPLIT distance="150" swimtime="00:02:01.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5921" number="1" />
                    <RELAYPOSITION athleteid="5884" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5879" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5898" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1368" points="302" swimtime="00:02:19.17" resultid="7434" heatid="10801" lane="0" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="150" swimtime="00:01:43.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5927" number="1" />
                    <RELAYPOSITION athleteid="5921" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5889" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5913" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" points="326" swimtime="00:02:03.25" resultid="7436" heatid="10871" lane="9" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                    <SPLIT distance="100" swimtime="00:00:57.45" />
                    <SPLIT distance="150" swimtime="00:01:31.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5927" number="1" />
                    <RELAYPOSITION athleteid="5921" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5889" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5913" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1518" points="212" swimtime="00:02:22.26" resultid="7433" heatid="10870" lane="7" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:13.09" />
                    <SPLIT distance="150" swimtime="00:01:48.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5905" number="1" />
                    <RELAYPOSITION athleteid="5884" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5879" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5898" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1347" points="141" swimtime="00:03:24.18" resultid="7429" heatid="10797" lane="4" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.13" />
                    <SPLIT distance="100" swimtime="00:01:40.08" />
                    <SPLIT distance="150" swimtime="00:02:20.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5846" number="1" />
                    <RELAYPOSITION athleteid="5831" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5837" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5826" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1497" points="421" swimtime="00:02:08.77" resultid="7435" heatid="10868" lane="0" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="100" swimtime="00:01:00.29" />
                    <SPLIT distance="150" swimtime="00:01:32.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5855" number="1" />
                    <RELAYPOSITION athleteid="5873" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5868" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5850" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1347" points="367" swimtime="00:02:28.50" resultid="7430" heatid="10798" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:21.85" />
                    <SPLIT distance="150" swimtime="00:01:53.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5855" number="1" />
                    <RELAYPOSITION athleteid="5868" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5873" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5850" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1497" points="123" swimtime="00:03:13.63" resultid="7432" heatid="10868" lane="4" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.57" />
                    <SPLIT distance="100" swimtime="00:01:31.55" />
                    <SPLIT distance="150" swimtime="00:02:09.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5846" number="1" />
                    <RELAYPOSITION athleteid="5831" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5837" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5826" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:20.48" resultid="7423" heatid="10732" lane="8" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:09.30" />
                    <SPLIT distance="150" swimtime="00:01:44.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5889" number="1" />
                    <RELAYPOSITION athleteid="5837" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5879" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5850" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1653" swimtime="00:02:46.58" resultid="7424" heatid="10928" lane="1" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.92" />
                    <SPLIT distance="150" swimtime="00:01:58.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5889" number="1" />
                    <RELAYPOSITION athleteid="5837" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5879" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5850" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:11.29" resultid="7425" heatid="10732" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:03.16" />
                    <SPLIT distance="150" swimtime="00:01:38.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5913" number="1" />
                    <RELAYPOSITION athleteid="5905" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5831" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5868" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1653" swimtime="00:02:50.76" resultid="7426" heatid="10928" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                    <SPLIT distance="100" swimtime="00:01:26.65" />
                    <SPLIT distance="150" swimtime="00:02:01.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5905" number="1" />
                    <RELAYPOSITION athleteid="5831" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5913" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5868" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:01:55.32" resultid="7427" heatid="10733" lane="6" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="100" swimtime="00:00:56.80" />
                    <SPLIT distance="150" swimtime="00:01:26.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5927" number="1" />
                    <RELAYPOSITION athleteid="5921" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5855" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5873" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1653" swimtime="00:02:15.72" resultid="7428" heatid="10929" lane="7" entrytime="00:02:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:10.69" />
                    <SPLIT distance="150" swimtime="00:01:43.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5927" number="1" />
                    <RELAYPOSITION athleteid="5921" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5855" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5873" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="RIKIP" nation="LAT" clubid="3785" name="Riga Kipsala Swimming Club">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Janis" gender="M" lastname="Plotnieks" nation="LAT" athleteid="3786">
              <RESULTS>
                <RESULT eventid="1190" points="391" swimtime="00:02:35.83" resultid="3787" heatid="10727" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="150" swimtime="00:01:57.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="418" swimtime="00:00:32.13" resultid="3788" heatid="10749" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1452" points="459" swimtime="00:01:07.21" resultid="3789" heatid="10850" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="369" swimtime="00:02:35.92" resultid="3790" heatid="10904" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:13.99" />
                    <SPLIT distance="150" swimtime="00:01:55.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RMRYB" nation="POL" region="SLA" clubid="3414" name="Rmks Rybnik">
          <CONTACT city="Rybnik" email="aniaduda0511@tlen.pl" name="Duda Anna" phone="792666159" state="SLA" street="orzepowicka 22a/37" zip="44-217" />
          <ATHLETES>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="3415">
              <RESULTS>
                <RESULT eventid="1144" points="571" swimtime="00:00:28.59" resultid="7961" heatid="10688" lane="2" entrytime="00:00:28.10" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat C  35-39  lat" eventid="1175" points="462" swimtime="00:02:43.08" resultid="7962" heatid="10718" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:15.02" />
                    <SPLIT distance="150" swimtime="00:02:05.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="420" swimtime="00:00:36.12" resultid="7963" heatid="10738" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1287" points="519" swimtime="00:01:04.75" resultid="7964" heatid="10771" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="548" swimtime="00:00:29.85" resultid="7965" heatid="10824" lane="4" entrytime="00:00:29.87" />
                <RESULT eventid="1437" points="396" swimtime="00:01:19.11" resultid="7966" heatid="10842" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="494" swimtime="00:01:10.16" resultid="7967" heatid="10884" lane="4" entrytime="00:01:09.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="454" swimtime="00:00:38.33" resultid="7968" heatid="10911" lane="1" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RYSEN" nation="POL" region="SLA" clubid="2982" name="Rydułtowska Akademia Aktywnego Seniora" shortname="Rydułtowska Akademia Aktywnego">
          <CONTACT email="otelom.080966@interia.pl" name="OTLIK MARIAN" />
          <ATHLETES>
            <ATHLETE birthdate="1946-02-02" firstname="Maria" gender="F" lastname="Lippa" nation="POL" athleteid="2993">
              <RESULTS>
                <RESULT eventid="1059" points="40" swimtime="00:23:32.53" resultid="7979" heatid="10665" lane="4" entrytime="00:21:10.00" />
                <RESULT eventid="1287" points="25" swimtime="00:02:55.86" resultid="7980" heatid="10765" lane="3" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="28" swimtime="00:03:11.00" resultid="7981" heatid="10839" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="35" swimtime="00:05:45.19" resultid="7982" heatid="10851" lane="7" entrytime="00:05:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.62" />
                    <SPLIT distance="100" swimtime="00:02:42.30" />
                    <SPLIT distance="150" swimtime="00:04:14.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="29" swimtime="00:06:42.93" resultid="7983" heatid="10893" lane="5" entrytime="00:06:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.50" />
                    <SPLIT distance="100" swimtime="00:03:18.88" />
                    <SPLIT distance="150" swimtime="00:05:05.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="38" swimtime="00:11:43.25" resultid="7984" heatid="10930" lane="4" entrytime="00:10:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.48" />
                    <SPLIT distance="100" swimtime="00:02:44.60" />
                    <SPLIT distance="150" swimtime="00:04:14.22" />
                    <SPLIT distance="200" swimtime="00:05:44.89" />
                    <SPLIT distance="250" swimtime="00:07:14.15" />
                    <SPLIT distance="300" swimtime="00:08:44.30" />
                    <SPLIT distance="350" swimtime="00:10:15.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-16" firstname="Bugla" gender="M" lastname="Rudolf" nation="POL" athleteid="2983">
              <RESULTS>
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="7970" heatid="10669" lane="7" entrytime="00:19:44.00" />
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="7971" heatid="10691" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1190" points="58" swimtime="00:04:53.86" resultid="7972" heatid="10720" lane="9" entrytime="00:04:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.41" />
                    <SPLIT distance="100" swimtime="00:02:30.74" />
                    <SPLIT distance="150" swimtime="00:03:51.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="73" swimtime="00:00:57.35" resultid="7973" heatid="10741" lane="7" entrytime="00:00:59.00" />
                <RESULT eventid="1332" status="DNS" swimtime="00:00:00.00" resultid="7974" heatid="10792" lane="0" entrytime="00:04:55.00" />
                <RESULT eventid="1422" points="53" swimtime="00:00:59.58" resultid="7975" heatid="10826" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1546" points="55" swimtime="00:10:40.70" resultid="7976" heatid="10876" lane="3" entrytime="00:09:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.44" />
                    <SPLIT distance="100" swimtime="00:02:37.21" />
                    <SPLIT distance="150" swimtime="00:04:03.78" />
                    <SPLIT distance="200" swimtime="00:05:29.19" />
                    <SPLIT distance="250" swimtime="00:06:53.25" />
                    <SPLIT distance="300" swimtime="00:08:16.30" />
                    <SPLIT distance="350" swimtime="00:09:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="32" swimtime="00:02:35.61" resultid="7977" heatid="10885" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="63" swimtime="00:04:39.92" resultid="7978" heatid="10899" lane="5" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.38" />
                    <SPLIT distance="100" swimtime="00:02:18.54" />
                    <SPLIT distance="150" swimtime="00:03:30.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-12-07" firstname="Miron" gender="M" lastname="Starosta" nation="POL" athleteid="3000">
              <RESULTS>
                <RESULT eventid="1160" points="83" swimtime="00:00:47.75" resultid="7985" heatid="10691" lane="8" entrytime="00:00:47.00" />
                <RESULT eventid="1190" points="62" swimtime="00:04:46.67" resultid="7986" heatid="10719" lane="5" entrytime="00:04:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.96" />
                    <SPLIT distance="100" swimtime="00:02:20.24" />
                    <SPLIT distance="150" swimtime="00:03:42.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="75" swimtime="00:04:59.85" resultid="7987" heatid="10757" lane="5" entrytime="00:04:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.46" />
                    <SPLIT distance="100" swimtime="00:02:20.82" />
                    <SPLIT distance="150" swimtime="00:03:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="72" swimtime="00:01:52.74" resultid="7988" heatid="10773" lane="6" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="71" swimtime="00:02:17.54" resultid="7989" heatid="10809" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="53" swimtime="00:10:47.59" resultid="7990" heatid="10876" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.70" />
                    <SPLIT distance="100" swimtime="00:02:41.74" />
                    <SPLIT distance="150" swimtime="00:04:11.50" />
                    <SPLIT distance="200" swimtime="00:05:36.82" />
                    <SPLIT distance="250" swimtime="00:07:03.82" />
                    <SPLIT distance="300" swimtime="00:08:27.78" />
                    <SPLIT distance="350" swimtime="00:09:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNF" swimtime="00:00:00.00" resultid="7991" heatid="10885" lane="8" />
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="7992" heatid="10899" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-23" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="3009">
              <RESULTS>
                <RESULT eventid="1098" points="180" swimtime="00:13:19.51" resultid="7993" heatid="10670" lane="3" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                    <SPLIT distance="100" swimtime="00:01:28.89" />
                    <SPLIT distance="150" swimtime="00:02:17.98" />
                    <SPLIT distance="200" swimtime="00:03:08.35" />
                    <SPLIT distance="250" swimtime="00:03:59.24" />
                    <SPLIT distance="300" swimtime="00:04:50.96" />
                    <SPLIT distance="350" swimtime="00:05:42.16" />
                    <SPLIT distance="400" swimtime="00:06:34.32" />
                    <SPLIT distance="450" swimtime="00:07:25.98" />
                    <SPLIT distance="500" swimtime="00:08:17.14" />
                    <SPLIT distance="550" swimtime="00:09:08.18" />
                    <SPLIT distance="600" swimtime="00:09:59.67" />
                    <SPLIT distance="650" swimtime="00:10:50.98" />
                    <SPLIT distance="700" swimtime="00:11:41.98" />
                    <SPLIT distance="750" swimtime="00:12:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="144" swimtime="00:03:37.43" resultid="7994" heatid="10722" lane="0" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                    <SPLIT distance="100" swimtime="00:01:41.24" />
                    <SPLIT distance="150" swimtime="00:02:47.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="165" swimtime="00:00:43.75" resultid="7995" heatid="10744" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1332" status="DNS" swimtime="00:00:00.00" resultid="7996" heatid="10792" lane="5" entrytime="00:03:55.00" />
                <RESULT eventid="1452" points="155" swimtime="00:01:36.43" resultid="7997" heatid="10846" lane="9" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" status="DNS" swimtime="00:00:00.00" resultid="7998" heatid="10877" lane="2" entrytime="00:07:21.00" />
                <RESULT eventid="1608" points="149" swimtime="00:03:31.06" resultid="7999" heatid="10901" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.11" />
                    <SPLIT distance="100" swimtime="00:01:43.13" />
                    <SPLIT distance="150" swimtime="00:02:38.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="8000" heatid="10939" lane="2" entrytime="00:06:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="6052" name="SC Marlin">
          <CONTACT city="Kyiv" email="kovalyovleonid@gmail.com, marlinsportclub@gmail.co" internet="www.marlinsc.com" name="Kovalyov Leonid" phone="+38 097 904 0114" street="79, Victory Avenue, Apt 48" zip="03000" />
          <ATHLETES>
            <ATHLETE birthdate="1986-12-24" firstname="Viktor" gender="M" lastname="Kucheriavyi" nation="UKR" athleteid="6053">
              <RESULTS>
                <RESULT eventid="1098" points="157" swimtime="00:13:56.92" resultid="6054" heatid="10670" lane="9" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:01:27.19" />
                    <SPLIT distance="150" swimtime="00:02:17.54" />
                    <SPLIT distance="200" swimtime="00:03:10.44" />
                    <SPLIT distance="250" swimtime="00:04:04.91" />
                    <SPLIT distance="300" swimtime="00:04:58.84" />
                    <SPLIT distance="350" swimtime="00:05:54.88" />
                    <SPLIT distance="400" swimtime="00:06:48.20" />
                    <SPLIT distance="450" swimtime="00:07:44.84" />
                    <SPLIT distance="500" swimtime="00:08:37.89" />
                    <SPLIT distance="550" swimtime="00:09:33.61" />
                    <SPLIT distance="600" swimtime="00:10:28.92" />
                    <SPLIT distance="650" swimtime="00:11:21.64" />
                    <SPLIT distance="700" swimtime="00:12:14.40" />
                    <SPLIT distance="750" swimtime="00:13:07.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="167" swimtime="00:00:43.65" resultid="6055" heatid="10744" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1302" points="243" swimtime="00:01:15.11" resultid="6056" heatid="10777" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="157" swimtime="00:01:36.07" resultid="6057" heatid="10845" lane="7" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="189" swimtime="00:02:57.67" resultid="6058" heatid="10859" lane="8" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                    <SPLIT distance="150" swimtime="00:02:12.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="150" swimtime="00:03:30.45" resultid="6059" heatid="10901" lane="9" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.41" />
                    <SPLIT distance="100" swimtime="00:01:41.44" />
                    <SPLIT distance="150" swimtime="00:02:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="169" swimtime="00:06:37.36" resultid="6060" heatid="10938" lane="7" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:27.84" />
                    <SPLIT distance="150" swimtime="00:02:18.39" />
                    <SPLIT distance="200" swimtime="00:03:10.81" />
                    <SPLIT distance="250" swimtime="00:04:04.78" />
                    <SPLIT distance="300" swimtime="00:04:58.17" />
                    <SPLIT distance="350" swimtime="00:05:50.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIGLI" nation="POL" region="SLA" clubid="3110" name="Sikret Gliwice">
          <CONTACT city="GLIWICE" email="JOANNAECO@TLEN.PL" internet="WWW.SIKRET-PLYWANIE.PL" name="ZAGAŁA JOANNA" phone="601427257" state="ŚLĄSK" street="JAGIELOŃSKA 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1981-02-14" firstname="Dawid" gender="M" lastname="Zimkowski" nation="POL" athleteid="3142">
              <RESULTS>
                <RESULT eventid="1190" points="267" swimtime="00:02:56.85" resultid="6508" heatid="10723" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:19.81" />
                    <SPLIT distance="150" swimtime="00:02:14.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="287" swimtime="00:00:36.44" resultid="6509" heatid="10748" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="273" swimtime="00:01:12.25" resultid="6510" heatid="10779" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="395" swimtime="00:00:30.57" resultid="6511" heatid="10831" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1452" points="237" swimtime="00:01:23.78" resultid="6512" heatid="10847" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="287" swimtime="00:05:33.43" resultid="6513" heatid="10941" lane="8" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:01:15.65" />
                    <SPLIT distance="150" swimtime="00:01:58.08" />
                    <SPLIT distance="200" swimtime="00:02:40.52" />
                    <SPLIT distance="250" swimtime="00:03:24.03" />
                    <SPLIT distance="300" swimtime="00:04:07.76" />
                    <SPLIT distance="350" swimtime="00:04:51.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-11" firstname="Agnieszka" gender="F" lastname="Drejka" nation="POL" athleteid="3128">
              <RESULTS>
                <RESULT eventid="1257" points="182" swimtime="00:04:05.40" resultid="6496" heatid="10754" lane="7" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.13" />
                    <SPLIT distance="100" swimtime="00:01:58.56" />
                    <SPLIT distance="150" swimtime="00:03:02.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="191" swimtime="00:01:30.39" resultid="6497" heatid="10766" lane="4" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="171" swimtime="00:01:55.83" resultid="6498" heatid="10804" lane="3" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="186" swimtime="00:03:17.63" resultid="6499" heatid="10852" lane="2" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                    <SPLIT distance="100" swimtime="00:01:31.88" />
                    <SPLIT distance="150" swimtime="00:02:25.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="168" swimtime="00:00:53.37" resultid="6500" heatid="10907" lane="8" entrytime="00:00:52.00" />
                <RESULT eventid="1674" points="165" swimtime="00:07:11.02" resultid="6501" heatid="10931" lane="2" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                    <SPLIT distance="100" swimtime="00:01:39.30" />
                    <SPLIT distance="150" swimtime="00:02:34.03" />
                    <SPLIT distance="200" swimtime="00:03:30.50" />
                    <SPLIT distance="250" swimtime="00:04:27.08" />
                    <SPLIT distance="300" swimtime="00:05:24.10" />
                    <SPLIT distance="350" swimtime="00:06:18.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-16" firstname="Stanisław" gender="M" lastname="Twardysko" nation="POL" athleteid="3135">
              <RESULTS>
                <RESULT eventid="1160" points="201" swimtime="00:00:35.68" resultid="6502" heatid="10695" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1242" points="118" swimtime="00:00:48.99" resultid="6503" heatid="10743" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1302" points="201" swimtime="00:01:19.99" resultid="6504" heatid="10776" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="153" swimtime="00:01:36.76" resultid="6505" heatid="10845" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="180" swimtime="00:03:00.41" resultid="6506" heatid="10858" lane="7" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                    <SPLIT distance="150" swimtime="00:02:13.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="137" swimtime="00:03:36.90" resultid="6507" heatid="10900" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.19" />
                    <SPLIT distance="150" swimtime="00:02:43.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="3111">
              <RESULTS>
                <RESULT eventid="1113" points="187" swimtime="00:26:55.62" resultid="6481" heatid="10674" lane="8" entrytime="00:30:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                    <SPLIT distance="100" swimtime="00:01:40.00" />
                    <SPLIT distance="150" swimtime="00:02:34.41" />
                    <SPLIT distance="200" swimtime="00:03:28.28" />
                    <SPLIT distance="250" swimtime="00:04:23.41" />
                    <SPLIT distance="300" swimtime="00:05:18.08" />
                    <SPLIT distance="350" swimtime="00:06:13.70" />
                    <SPLIT distance="400" swimtime="00:07:08.71" />
                    <SPLIT distance="450" swimtime="00:08:04.58" />
                    <SPLIT distance="500" swimtime="00:08:59.91" />
                    <SPLIT distance="550" swimtime="00:09:54.64" />
                    <SPLIT distance="600" swimtime="00:10:49.28" />
                    <SPLIT distance="650" swimtime="00:11:43.92" />
                    <SPLIT distance="700" swimtime="00:12:38.71" />
                    <SPLIT distance="750" swimtime="00:13:33.90" />
                    <SPLIT distance="800" swimtime="00:14:28.38" />
                    <SPLIT distance="850" swimtime="00:15:22.93" />
                    <SPLIT distance="900" swimtime="00:16:16.92" />
                    <SPLIT distance="950" swimtime="00:17:11.17" />
                    <SPLIT distance="1000" swimtime="00:18:05.43" />
                    <SPLIT distance="1050" swimtime="00:18:58.78" />
                    <SPLIT distance="1100" swimtime="00:19:52.42" />
                    <SPLIT distance="1150" swimtime="00:20:46.84" />
                    <SPLIT distance="1200" swimtime="00:21:40.46" />
                    <SPLIT distance="1250" swimtime="00:22:33.85" />
                    <SPLIT distance="1300" swimtime="00:23:27.26" />
                    <SPLIT distance="1350" swimtime="00:24:21.38" />
                    <SPLIT distance="1400" swimtime="00:25:14.42" />
                    <SPLIT distance="1450" swimtime="00:26:07.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="216" swimtime="00:00:39.52" resultid="6482" heatid="10683" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1226" points="172" swimtime="00:00:48.65" resultid="6483" heatid="10734" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1287" points="224" swimtime="00:01:25.70" resultid="6484" heatid="10767" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="164" swimtime="00:01:46.05" resultid="6485" heatid="10839" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="201" swimtime="00:03:12.81" resultid="6486" heatid="10852" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                    <SPLIT distance="100" swimtime="00:01:35.64" />
                    <SPLIT distance="150" swimtime="00:02:27.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="158" swimtime="00:03:49.13" resultid="6487" heatid="10894" lane="4" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.08" />
                    <SPLIT distance="100" swimtime="00:01:56.13" />
                    <SPLIT distance="150" swimtime="00:02:54.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="193" swimtime="00:00:50.99" resultid="6488" heatid="10906" lane="7" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="3120">
              <RESULTS>
                <RESULT eventid="1144" points="174" swimtime="00:00:42.49" resultid="6489" heatid="10683" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="1257" points="152" swimtime="00:04:20.64" resultid="6490" heatid="10753" lane="3" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.88" />
                    <SPLIT distance="100" swimtime="00:02:08.69" />
                    <SPLIT distance="150" swimtime="00:03:14.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1317" status="DNS" swimtime="00:00:00.00" resultid="6491" heatid="10789" lane="5" entrytime="00:05:00.00" />
                <RESULT eventid="1376" points="151" swimtime="00:02:00.82" resultid="6492" heatid="10804" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="90" swimtime="00:09:54.15" resultid="6493" heatid="10873" lane="3" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.66" />
                    <SPLIT distance="100" swimtime="00:02:29.40" />
                    <SPLIT distance="150" swimtime="00:03:58.17" />
                    <SPLIT distance="200" swimtime="00:05:27.47" />
                    <SPLIT distance="250" swimtime="00:06:37.90" />
                    <SPLIT distance="300" swimtime="00:07:48.15" />
                    <SPLIT distance="350" swimtime="00:08:53.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="69" swimtime="00:02:14.73" resultid="6494" heatid="10883" lane="9" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="185" swimtime="00:00:51.66" resultid="6495" heatid="10907" lane="7" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:27.17" resultid="6514" heatid="10731" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.38" />
                    <SPLIT distance="150" swimtime="00:01:56.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3120" number="1" />
                    <RELAYPOSITION athleteid="3135" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3111" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3142" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1653" swimtime="00:02:50.89" resultid="6515" heatid="10928" lane="9" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.11" />
                    <SPLIT distance="100" swimtime="00:01:43.86" />
                    <SPLIT distance="150" swimtime="00:02:14.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3111" number="1" />
                    <RELAYPOSITION athleteid="3120" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3142" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3135" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="STEEF" nation="POL" region="DOL" clubid="4592" name="Steef">
          <CONTACT city="Wrocław" email="ste1@wp.pl" name="Stefan Skrzypek" street="Edyty Stein 6/1" zip="50-322" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="4600">
              <RESULTS>
                <RESULT eventid="1128" points="162" swimtime="00:26:37.02" resultid="8093" heatid="10676" lane="6" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.07" />
                    <SPLIT distance="100" swimtime="00:01:36.42" />
                    <SPLIT distance="150" swimtime="00:02:28.14" />
                    <SPLIT distance="200" swimtime="00:03:19.97" />
                    <SPLIT distance="250" swimtime="00:04:11.15" />
                    <SPLIT distance="300" swimtime="00:05:04.07" />
                    <SPLIT distance="350" swimtime="00:05:57.36" />
                    <SPLIT distance="400" swimtime="00:06:50.48" />
                    <SPLIT distance="450" swimtime="00:07:45.60" />
                    <SPLIT distance="500" swimtime="00:08:38.57" />
                    <SPLIT distance="550" swimtime="00:09:33.27" />
                    <SPLIT distance="600" swimtime="00:10:26.59" />
                    <SPLIT distance="650" swimtime="00:11:20.42" />
                    <SPLIT distance="700" swimtime="00:12:13.02" />
                    <SPLIT distance="750" swimtime="00:13:07.69" />
                    <SPLIT distance="800" swimtime="00:14:01.59" />
                    <SPLIT distance="850" swimtime="00:14:54.94" />
                    <SPLIT distance="900" swimtime="00:15:49.72" />
                    <SPLIT distance="950" swimtime="00:16:48.07" />
                    <SPLIT distance="1000" swimtime="00:17:42.56" />
                    <SPLIT distance="1050" swimtime="00:18:35.68" />
                    <SPLIT distance="1100" swimtime="00:19:28.64" />
                    <SPLIT distance="1150" swimtime="00:20:22.94" />
                    <SPLIT distance="1200" swimtime="00:21:16.07" />
                    <SPLIT distance="1250" swimtime="00:22:10.00" />
                    <SPLIT distance="1300" swimtime="00:23:04.19" />
                    <SPLIT distance="1350" swimtime="00:23:58.58" />
                    <SPLIT distance="1400" swimtime="00:24:53.47" />
                    <SPLIT distance="1450" swimtime="00:25:46.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="8094" heatid="10758" lane="6" entrytime="00:03:50.00" />
                <RESULT eventid="1482" points="177" swimtime="00:03:01.40" resultid="8095" heatid="10858" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                    <SPLIT distance="100" swimtime="00:01:28.13" />
                    <SPLIT distance="150" swimtime="00:02:14.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="8096" heatid="10914" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="1695" points="162" swimtime="00:06:43.02" resultid="8097" heatid="10938" lane="8" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                    <SPLIT distance="100" swimtime="00:01:36.78" />
                    <SPLIT distance="150" swimtime="00:02:28.47" />
                    <SPLIT distance="200" swimtime="00:03:22.37" />
                    <SPLIT distance="250" swimtime="00:04:13.96" />
                    <SPLIT distance="300" swimtime="00:05:06.34" />
                    <SPLIT distance="350" swimtime="00:05:55.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="4593">
              <RESULTS>
                <RESULT eventid="1175" points="305" swimtime="00:03:07.19" resultid="8087" heatid="10716" lane="1" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                    <SPLIT distance="100" swimtime="00:01:28.02" />
                    <SPLIT distance="150" swimtime="00:02:22.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="298" swimtime="00:00:40.48" resultid="8088" heatid="10736" lane="4" entrytime="00:00:42.50" />
                <RESULT eventid="1437" points="295" swimtime="00:01:27.29" resultid="8089" heatid="10841" lane="2" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="274" swimtime="00:06:49.72" resultid="8090" heatid="10874" lane="3" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                    <SPLIT distance="100" swimtime="00:01:36.67" />
                    <SPLIT distance="150" swimtime="00:02:27.42" />
                    <SPLIT distance="200" swimtime="00:03:17.11" />
                    <SPLIT distance="250" swimtime="00:04:14.90" />
                    <SPLIT distance="300" swimtime="00:05:13.33" />
                    <SPLIT distance="350" swimtime="00:06:02.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="280" swimtime="00:03:09.56" resultid="8091" heatid="10896" lane="2" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                    <SPLIT distance="100" swimtime="00:01:30.84" />
                    <SPLIT distance="150" swimtime="00:02:20.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="254" swimtime="00:06:13.26" resultid="8092" heatid="10932" lane="6" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                    <SPLIT distance="100" swimtime="00:01:30.63" />
                    <SPLIT distance="150" swimtime="00:02:18.70" />
                    <SPLIT distance="200" swimtime="00:03:06.92" />
                    <SPLIT distance="250" swimtime="00:03:55.19" />
                    <SPLIT distance="300" swimtime="00:04:41.82" />
                    <SPLIT distance="350" swimtime="00:05:27.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SMMK" nation="POL" region="KR" clubid="4269" name="Straż Miejska Miasta Kraków">
          <CONTACT city="Kraków" name="Jawień Krzysztof" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1971-06-11" firstname="Krzysztof" gender="M" lastname="Jawień" nation="POL" athleteid="4285">
              <RESULTS>
                <RESULT eventid="1098" points="250" swimtime="00:11:57.20" resultid="6738" heatid="10670" lane="1" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                    <SPLIT distance="150" swimtime="00:01:59.56" />
                    <SPLIT distance="200" swimtime="00:02:44.03" />
                    <SPLIT distance="250" swimtime="00:03:28.84" />
                    <SPLIT distance="300" swimtime="00:04:14.17" />
                    <SPLIT distance="350" swimtime="00:04:59.03" />
                    <SPLIT distance="400" swimtime="00:05:44.56" />
                    <SPLIT distance="450" swimtime="00:06:30.14" />
                    <SPLIT distance="500" swimtime="00:07:16.43" />
                    <SPLIT distance="550" swimtime="00:08:02.65" />
                    <SPLIT distance="600" swimtime="00:08:49.90" />
                    <SPLIT distance="650" swimtime="00:09:37.85" />
                    <SPLIT distance="700" swimtime="00:10:25.98" />
                    <SPLIT distance="750" swimtime="00:11:12.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="305" swimtime="00:02:49.22" resultid="6739" heatid="10724" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:19.31" />
                    <SPLIT distance="150" swimtime="00:02:08.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="317" swimtime="00:03:06.15" resultid="6740" heatid="10757" lane="4" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:29.75" />
                    <SPLIT distance="150" swimtime="00:02:18.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="201" swimtime="00:03:10.36" resultid="6741" heatid="10794" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="100" swimtime="00:01:24.28" />
                    <SPLIT distance="150" swimtime="00:02:16.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="316" swimtime="00:01:23.84" resultid="6742" heatid="10816" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="292" swimtime="00:06:07.28" resultid="6743" heatid="10879" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                    <SPLIT distance="150" swimtime="00:02:09.24" />
                    <SPLIT distance="200" swimtime="00:02:59.24" />
                    <SPLIT distance="250" swimtime="00:03:49.27" />
                    <SPLIT distance="300" swimtime="00:04:40.24" />
                    <SPLIT distance="350" swimtime="00:05:23.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="255" swimtime="00:02:56.48" resultid="6744" heatid="10900" lane="9" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:23.30" />
                    <SPLIT distance="150" swimtime="00:02:10.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="337" swimtime="00:00:37.93" resultid="6745" heatid="10922" lane="8" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STSWI" nation="POL" region="14" clubid="9227" name="Swimmers St Pływackie">
          <CONTACT city="WARSZAWA" email="REMOG@SWIMMERSTEAM.PL" name="GOŁĘBIOWSKI REMO" phone="601333782" state="MAZ" street="GŁADKA 18" zip="02-172" />
          <ATHLETES>
            <ATHLETE birthdate="1982-07-12" firstname="Katarzyna" gender="M" lastname="Hereczyńska" nation="POL" athleteid="9455">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="9456" heatid="10695" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-12" firstname="Jan" gender="M" lastname="Rekowski" nation="POL" athleteid="9432">
              <RESULTS>
                <RESULT eventid="1160" points="471" swimtime="00:00:26.86" resultid="9433" heatid="10709" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1190" points="311" swimtime="00:02:48.12" resultid="9434" heatid="10726" lane="0" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:16.81" />
                    <SPLIT distance="150" swimtime="00:02:07.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="351" swimtime="00:00:34.05" resultid="9435" heatid="10747" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="466" swimtime="00:01:00.49" resultid="9436" heatid="10785" lane="5" entrytime="00:00:59.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-10-21" firstname="Piotr" gender="M" lastname="Macioszek" nation="POL" athleteid="9403">
              <RESULTS>
                <RESULT eventid="1160" points="176" swimtime="00:00:37.25" resultid="9404" heatid="10696" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1190" points="118" swimtime="00:03:51.91" resultid="9405" heatid="10723" lane="7" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.93" />
                    <SPLIT distance="100" swimtime="00:01:52.62" />
                    <SPLIT distance="150" swimtime="00:02:56.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="97" swimtime="00:00:52.32" resultid="9406" heatid="10745" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="1392" points="141" swimtime="00:01:49.63" resultid="9407" heatid="10813" lane="9" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="95" swimtime="00:01:53.54" resultid="9408" heatid="10846" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="163" swimtime="00:00:48.28" resultid="9409" heatid="10916" lane="8" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Marek" gender="M" lastname="Brożyna" nation="POL" athleteid="9426">
              <RESULTS>
                <RESULT eventid="1190" points="316" swimtime="00:02:47.32" resultid="9427" heatid="10726" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:16.63" />
                    <SPLIT distance="150" swimtime="00:02:09.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="341" swimtime="00:00:34.38" resultid="9428" heatid="10748" lane="1" entrytime="00:00:34.30" />
                <RESULT eventid="1452" points="343" swimtime="00:01:14.07" resultid="9429" heatid="10848" lane="9" entrytime="00:01:16.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="294" swimtime="00:06:06.33" resultid="9430" heatid="10876" lane="1">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:11.33" />
                    <SPLIT distance="200" swimtime="00:02:56.52" />
                    <SPLIT distance="250" swimtime="00:03:51.36" />
                    <SPLIT distance="300" swimtime="00:04:46.08" />
                    <SPLIT distance="350" swimtime="00:05:26.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="340" swimtime="00:02:40.24" resultid="9431" heatid="10903" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                    <SPLIT distance="100" swimtime="00:01:18.68" />
                    <SPLIT distance="150" swimtime="00:02:00.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="Piotr" gender="M" lastname="Gajewski" nation="POL" athleteid="9512">
              <RESULTS>
                <RESULT eventid="1128" points="276" swimtime="00:22:17.06" resultid="9513" heatid="10678" lane="7" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:25.34" />
                    <SPLIT distance="150" swimtime="00:02:09.48" />
                    <SPLIT distance="200" swimtime="00:02:54.41" />
                    <SPLIT distance="250" swimtime="00:03:39.21" />
                    <SPLIT distance="300" swimtime="00:04:24.02" />
                    <SPLIT distance="350" swimtime="00:05:09.00" />
                    <SPLIT distance="400" swimtime="00:05:54.08" />
                    <SPLIT distance="450" swimtime="00:06:39.29" />
                    <SPLIT distance="500" swimtime="00:07:24.65" />
                    <SPLIT distance="550" swimtime="00:08:09.94" />
                    <SPLIT distance="600" swimtime="00:08:55.24" />
                    <SPLIT distance="650" swimtime="00:09:40.69" />
                    <SPLIT distance="700" swimtime="00:10:26.30" />
                    <SPLIT distance="750" swimtime="00:11:11.72" />
                    <SPLIT distance="800" swimtime="00:11:57.29" />
                    <SPLIT distance="850" swimtime="00:12:42.08" />
                    <SPLIT distance="900" swimtime="00:13:27.33" />
                    <SPLIT distance="950" swimtime="00:14:11.38" />
                    <SPLIT distance="1000" swimtime="00:14:55.97" />
                    <SPLIT distance="1050" swimtime="00:15:40.38" />
                    <SPLIT distance="1100" swimtime="00:16:25.08" />
                    <SPLIT distance="1150" swimtime="00:17:09.39" />
                    <SPLIT distance="1200" swimtime="00:17:54.34" />
                    <SPLIT distance="1250" swimtime="00:18:38.38" />
                    <SPLIT distance="1300" swimtime="00:19:22.52" />
                    <SPLIT distance="1350" swimtime="00:20:06.60" />
                    <SPLIT distance="1400" swimtime="00:20:50.81" />
                    <SPLIT distance="1450" swimtime="00:21:34.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="324" swimtime="00:02:42.81" resultid="9514" heatid="10903" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:19.38" />
                    <SPLIT distance="150" swimtime="00:02:01.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="362" swimtime="00:01:12.74" resultid="9515" heatid="10848" lane="6" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-19" firstname="Krzysztof" gender="M" lastname="Jarocki" nation="POL" athleteid="9415">
              <RESULTS>
                <RESULT eventid="1160" points="107" swimtime="00:00:43.95" resultid="9416" heatid="10692" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="9417" heatid="10743" lane="3" entrytime="00:00:44.00" />
                <RESULT eventid="1638" points="120" swimtime="00:00:53.49" resultid="9418" heatid="10915" lane="9" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-27" firstname="Remigiusz" gender="M" lastname="Miklewski" nation="POL" athleteid="9398">
              <RESULTS>
                <RESULT eventid="1160" points="327" swimtime="00:00:30.33" resultid="9399" heatid="10701" lane="7" entrytime="00:00:29.90" />
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="9400" heatid="10747" lane="1" entrytime="00:00:35.90" />
                <RESULT eventid="1422" points="249" swimtime="00:00:35.61" resultid="9401" heatid="10829" lane="4" entrytime="00:00:34.90" />
                <RESULT eventid="1638" points="256" swimtime="00:00:41.57" resultid="9402" heatid="10918" lane="4" entrytime="00:00:39.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Arkadiusz" gender="M" lastname="Aptewicz" nation="POL" athleteid="9517">
              <RESULTS>
                <RESULT eventid="1190" points="534" swimtime="00:02:20.51" resultid="9518" heatid="10730" lane="4" entrytime="00:02:17.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                    <SPLIT distance="100" swimtime="00:01:07.14" />
                    <SPLIT distance="150" swimtime="00:01:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="580" swimtime="00:02:32.24" resultid="9519" heatid="10764" lane="5" entrytime="00:02:27.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:51.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="518" swimtime="00:01:11.09" resultid="9520" heatid="10819" lane="6" entrytime="00:01:09.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="543" swimtime="00:04:58.73" resultid="9521" heatid="10881" lane="5" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:07.44" />
                    <SPLIT distance="150" swimtime="00:01:50.67" />
                    <SPLIT distance="200" swimtime="00:02:32.93" />
                    <SPLIT distance="250" swimtime="00:03:12.13" />
                    <SPLIT distance="300" swimtime="00:03:52.55" />
                    <SPLIT distance="350" swimtime="00:04:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="583" swimtime="00:04:23.31" resultid="9522" heatid="10945" lane="4" entrytime="00:04:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                    <SPLIT distance="100" swimtime="00:01:04.73" />
                    <SPLIT distance="150" swimtime="00:01:38.30" />
                    <SPLIT distance="200" swimtime="00:02:11.76" />
                    <SPLIT distance="250" swimtime="00:02:44.74" />
                    <SPLIT distance="300" swimtime="00:03:18.07" />
                    <SPLIT distance="350" swimtime="00:03:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="541" swimtime="00:00:32.41" resultid="9523" heatid="10926" lane="7" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-10" firstname="Adam" gender="M" lastname="Komorowski" nation="POL" athleteid="9419">
              <RESULTS>
                <RESULT eventid="1128" points="120" swimtime="00:29:25.18" resultid="9420" heatid="10675" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:01:28.18" />
                    <SPLIT distance="150" swimtime="00:02:22.18" />
                    <SPLIT distance="200" swimtime="00:03:18.73" />
                    <SPLIT distance="250" swimtime="00:04:15.90" />
                    <SPLIT distance="300" swimtime="00:05:15.53" />
                    <SPLIT distance="350" swimtime="00:06:16.14" />
                    <SPLIT distance="400" swimtime="00:07:17.04" />
                    <SPLIT distance="450" swimtime="00:08:18.56" />
                    <SPLIT distance="500" swimtime="00:09:18.44" />
                    <SPLIT distance="550" swimtime="00:10:19.50" />
                    <SPLIT distance="600" swimtime="00:11:19.12" />
                    <SPLIT distance="650" swimtime="00:12:19.56" />
                    <SPLIT distance="700" swimtime="00:13:19.15" />
                    <SPLIT distance="750" swimtime="00:14:19.58" />
                    <SPLIT distance="800" swimtime="00:15:19.04" />
                    <SPLIT distance="850" swimtime="00:16:19.56" />
                    <SPLIT distance="900" swimtime="00:17:18.75" />
                    <SPLIT distance="950" swimtime="00:18:19.64" />
                    <SPLIT distance="1000" swimtime="00:19:20.45" />
                    <SPLIT distance="1050" swimtime="00:20:20.72" />
                    <SPLIT distance="1100" swimtime="00:21:20.41" />
                    <SPLIT distance="1150" swimtime="00:22:22.07" />
                    <SPLIT distance="1200" swimtime="00:23:22.54" />
                    <SPLIT distance="1250" swimtime="00:24:24.12" />
                    <SPLIT distance="1300" swimtime="00:25:24.18" />
                    <SPLIT distance="1350" swimtime="00:26:25.94" />
                    <SPLIT distance="1400" swimtime="00:27:26.42" />
                    <SPLIT distance="1450" swimtime="00:28:27.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="216" swimtime="00:00:34.82" resultid="9421" heatid="10697" lane="2" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-10" firstname="Małgorzata" gender="F" lastname="Cichocka" nation="POL" athleteid="9389">
              <RESULTS>
                <RESULT eventid="1144" points="289" swimtime="00:00:35.88" resultid="9390" heatid="10684" lane="0" entrytime="00:00:37.50" />
                <RESULT eventid="1226" points="228" swimtime="00:00:44.28" resultid="9391" heatid="10737" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1376" points="172" swimtime="00:01:55.64" resultid="9392" heatid="10806" lane="3" entrytime="00:01:35.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="9393" heatid="10908" lane="0" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-24" firstname="Katarzyna" gender="F" lastname="Bryłka" nation="POL" athleteid="9437">
              <RESULTS>
                <RESULT eventid="1144" points="93" swimtime="00:00:52.26" resultid="9438" heatid="10682" lane="3" entrytime="00:00:43.00" />
                <RESULT eventid="1226" points="108" swimtime="00:00:56.69" resultid="9439" heatid="10736" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1623" points="210" swimtime="00:00:49.56" resultid="9440" heatid="10907" lane="5" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-23" firstname="Justyna" gender="F" lastname="Sztuka-Wojtas" nation="POL" athleteid="9410">
              <RESULTS>
                <RESULT eventid="1144" points="234" swimtime="00:00:38.48" resultid="9411" heatid="10683" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="1287" points="198" swimtime="00:01:29.22" resultid="9412" heatid="10767" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="271" swimtime="00:01:39.35" resultid="9413" heatid="10806" lane="1" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="271" swimtime="00:00:45.54" resultid="9414" heatid="10908" lane="6" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-07-07" firstname="Remigiusz" gender="M" lastname="Gołębiowski" nation="POL" license="507914700017" athleteid="9380">
              <RESULTS>
                <RESULT eventid="1160" points="411" swimtime="00:00:28.12" resultid="9381" heatid="10705" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1302" points="434" swimtime="00:01:01.93" resultid="9382" heatid="10785" lane="1" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="458" swimtime="00:00:29.08" resultid="9383" heatid="10836" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1482" points="362" swimtime="00:02:23.11" resultid="9384" heatid="10865" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="100" swimtime="00:01:07.28" />
                    <SPLIT distance="150" swimtime="00:01:44.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-10-22" firstname="Katarzyna" gender="F" lastname="Frączyk" nation="POL" athleteid="9422">
              <RESULTS>
                <RESULT eventid="1144" points="261" swimtime="00:00:37.10" resultid="9423" heatid="10683" lane="0" entrytime="00:00:41.00" />
                <RESULT eventid="1407" points="116" swimtime="00:00:49.99" resultid="9424" heatid="10821" lane="2" entrytime="00:00:46.00" />
                <RESULT eventid="1467" points="140" swimtime="00:03:37.30" resultid="9425" heatid="10853" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.99" />
                    <SPLIT distance="100" swimtime="00:01:39.78" />
                    <SPLIT distance="150" swimtime="00:02:39.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-04" firstname="Norbert" gender="M" lastname="Tchorzewski" nation="POL" athleteid="9445">
              <RESULTS>
                <RESULT eventid="1128" points="195" swimtime="00:24:59.80" resultid="9446" heatid="10677" lane="1" entrytime="00:23:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:01:25.70" />
                    <SPLIT distance="150" swimtime="00:02:12.34" />
                    <SPLIT distance="200" swimtime="00:02:58.79" />
                    <SPLIT distance="250" swimtime="00:03:46.72" />
                    <SPLIT distance="300" swimtime="00:04:35.89" />
                    <SPLIT distance="350" swimtime="00:05:26.55" />
                    <SPLIT distance="400" swimtime="00:06:17.29" />
                    <SPLIT distance="450" swimtime="00:07:08.80" />
                    <SPLIT distance="500" swimtime="00:08:00.04" />
                    <SPLIT distance="550" swimtime="00:08:51.28" />
                    <SPLIT distance="600" swimtime="00:09:43.14" />
                    <SPLIT distance="650" swimtime="00:10:35.75" />
                    <SPLIT distance="700" swimtime="00:11:27.78" />
                    <SPLIT distance="750" swimtime="00:12:18.65" />
                    <SPLIT distance="800" swimtime="00:13:10.69" />
                    <SPLIT distance="850" swimtime="00:14:01.81" />
                    <SPLIT distance="900" swimtime="00:14:52.45" />
                    <SPLIT distance="950" swimtime="00:15:43.06" />
                    <SPLIT distance="1000" swimtime="00:16:33.38" />
                    <SPLIT distance="1050" swimtime="00:17:24.39" />
                    <SPLIT distance="1100" swimtime="00:18:15.05" />
                    <SPLIT distance="1150" swimtime="00:19:06.01" />
                    <SPLIT distance="1200" swimtime="00:19:58.23" />
                    <SPLIT distance="1250" swimtime="00:20:48.06" />
                    <SPLIT distance="1300" swimtime="00:21:39.64" />
                    <SPLIT distance="1350" swimtime="00:22:30.04" />
                    <SPLIT distance="1400" swimtime="00:23:20.83" />
                    <SPLIT distance="1450" swimtime="00:24:12.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="294" swimtime="00:00:31.44" resultid="9447" heatid="10701" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1190" points="191" swimtime="00:03:17.85" resultid="9448" heatid="10724" lane="9" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:31.92" />
                    <SPLIT distance="150" swimtime="00:02:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="9449" heatid="10780" lane="1" entrytime="00:01:07.90" />
                <RESULT eventid="1332" points="165" swimtime="00:03:23.24" resultid="9450" heatid="10793" lane="3" entrytime="00:03:14.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                    <SPLIT distance="100" swimtime="00:01:35.50" />
                    <SPLIT distance="150" swimtime="00:02:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="281" swimtime="00:00:34.23" resultid="9451" heatid="10828" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="9452" heatid="10861" lane="0" entrytime="00:02:38.00" />
                <RESULT eventid="1578" points="199" swimtime="00:01:25.23" resultid="9453" heatid="10888" lane="0" entrytime="00:01:19.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="9454" heatid="10941" lane="9" entrytime="00:05:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-03" firstname="Bolesław" gender="M" lastname="Porolniczak" nation="POL" athleteid="9394">
              <RESULTS>
                <RESULT eventid="1160" points="408" swimtime="00:00:28.18" resultid="9395" heatid="10707" lane="0" entrytime="00:00:27.30" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="9396" heatid="10783" lane="4" entrytime="00:01:02.78" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="9397" heatid="10833" lane="7" entrytime="00:00:30.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-09-14" firstname="Izabela" gender="F" lastname="Zyga" nation="POL" athleteid="9385">
              <RESULTS>
                <RESULT eventid="1257" points="469" swimtime="00:02:58.96" resultid="9386" heatid="10756" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:01:27.10" />
                    <SPLIT distance="150" swimtime="00:02:13.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="500" swimtime="00:01:21.04" resultid="9387" heatid="10808" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="451" swimtime="00:00:38.42" resultid="9388" heatid="10911" lane="5" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-12-11" firstname="Mikołaj" gender="M" lastname="Tusiński" nation="POL" athleteid="9441">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="9442" heatid="10700" lane="6" entrytime="00:00:30.30" />
                <RESULT eventid="1302" points="390" swimtime="00:01:04.16" resultid="9443" heatid="10783" lane="7" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="358" swimtime="00:00:31.58" resultid="9444" heatid="10831" lane="1" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" name="WARIATY 1" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="402" swimtime="00:02:06.51" resultid="9460" heatid="10799" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9426" number="1" />
                    <RELAYPOSITION athleteid="9432" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9380" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9441" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" points="400" swimtime="00:01:55.13" resultid="9461" heatid="10869" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                    <SPLIT distance="100" swimtime="00:00:56.72" />
                    <SPLIT distance="150" swimtime="00:01:25.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9380" number="1" />
                    <RELAYPOSITION athleteid="9441" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9426" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9512" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" name="WARIATY 2" number="2">
              <RESULTS>
                <RESULT eventid="1518" points="263" swimtime="00:02:12.39" resultid="9463" heatid="10869" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:03.95" />
                    <SPLIT distance="150" swimtime="00:01:42.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9445" number="1" />
                    <RELAYPOSITION athleteid="9419" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9403" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9398" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1347" status="DNS" swimtime="00:00:00.00" resultid="11200" heatid="10798" lane="0" late="yes">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9437" number="1" />
                    <RELAYPOSITION athleteid="9389" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9410" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9422" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" name="PANIE" number="1">
              <RESULTS>
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="9464" heatid="10867" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9437" number="1" />
                    <RELAYPOSITION athleteid="9422" number="2" />
                    <RELAYPOSITION athleteid="9389" number="3" />
                    <RELAYPOSITION athleteid="9410" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" name="PANIE 1" number="1">
              <RESULTS>
                <RESULT eventid="1347" points="189" status="EXH" swimtime="00:03:05.05" resultid="9459" heatid="10797" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.28" />
                    <SPLIT distance="100" swimtime="00:01:41.62" />
                    <SPLIT distance="150" swimtime="00:02:27.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9437" number="1" />
                    <RELAYPOSITION athleteid="9410" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9389" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9422" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="WARIAT 1" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:47.95" resultid="9457" heatid="10731" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.99" />
                    <SPLIT distance="100" swimtime="00:01:36.69" />
                    <SPLIT distance="150" swimtime="00:02:14.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9415" number="1" />
                    <RELAYPOSITION athleteid="9437" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9422" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9419" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="WARIATY 1" number="1">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:23.32" resultid="9465" heatid="10927" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.81" />
                    <SPLIT distance="150" swimtime="00:01:48.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9512" number="1" />
                    <RELAYPOSITION athleteid="9410" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9380" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9422" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="WARIAT 2" number="2">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="9458" heatid="10731" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9432" number="1" />
                    <RELAYPOSITION athleteid="9410" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9389" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9380" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="WARIATY 2" number="2">
              <RESULTS>
                <RESULT eventid="1653" status="DNS" swimtime="00:00:00.00" resultid="9466" heatid="10927" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9437" number="1" />
                    <RELAYPOSITION athleteid="9422" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="9445" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="9419" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SWSZC" nation="POL" region="ZAC" clubid="3819" name="Swimming Masters Team Szczecin">
          <CONTACT city="Szczecin" email="aga.krzyzostaniak@gmail.com" name="Krzyżostaniak Agnieszka" phone="603772862" street="Żupańskiego 12/8" zip="71-440" />
          <ATHLETES>
            <ATHLETE birthdate="1986-04-18" firstname="Jan" gender="M" lastname="Roenig" nation="POL" athleteid="3825">
              <RESULTS>
                <RESULT eventid="1160" points="426" swimtime="00:00:27.77" resultid="3826" heatid="10700" lane="2" entrytime="00:00:30.45" />
                <RESULT eventid="1302" points="389" swimtime="00:01:04.25" resultid="3827" heatid="10780" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="300" swimtime="00:01:25.33" resultid="3828" heatid="10813" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="430" swimtime="00:00:34.98" resultid="3829" heatid="10919" lane="6" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-12" firstname="Marek" gender="M" lastname="Zienkiewicz" nation="POL" athleteid="3852">
              <RESULTS>
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="3853" heatid="10670" lane="4" entrytime="00:12:00.00" />
                <RESULT eventid="1160" points="319" swimtime="00:00:30.59" resultid="3854" heatid="10700" lane="8" entrytime="00:00:30.58" />
                <RESULT eventid="1190" points="210" swimtime="00:03:11.78" resultid="3855" heatid="10722" lane="8" entrytime="00:03:12.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:29.79" />
                    <SPLIT distance="150" swimtime="00:02:22.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="289" swimtime="00:01:10.94" resultid="3856" heatid="10778" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="292" swimtime="00:00:33.80" resultid="3857" heatid="10830" lane="9" entrytime="00:00:34.90" />
                <RESULT eventid="1482" points="224" swimtime="00:02:47.84" resultid="3858" heatid="10859" lane="5" entrytime="00:02:50.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:17.11" />
                    <SPLIT distance="150" swimtime="00:02:01.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="312" swimtime="00:00:38.94" resultid="3859" heatid="10917" lane="4" entrytime="00:00:40.06" />
                <RESULT eventid="1695" points="206" swimtime="00:06:12.62" resultid="3860" heatid="10939" lane="3" entrytime="00:06:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:21.89" />
                    <SPLIT distance="150" swimtime="00:02:07.76" />
                    <SPLIT distance="200" swimtime="00:02:55.05" />
                    <SPLIT distance="250" swimtime="00:03:42.94" />
                    <SPLIT distance="300" swimtime="00:04:32.83" />
                    <SPLIT distance="350" swimtime="00:05:23.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-29" firstname="Robert" gender="M" lastname="Szota" nation="POL" athleteid="3836">
              <RESULTS>
                <RESULT eventid="1098" points="332" swimtime="00:10:52.51" resultid="3837" heatid="10671" lane="2" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:01:56.43" />
                    <SPLIT distance="200" swimtime="00:02:38.56" />
                    <SPLIT distance="250" swimtime="00:03:20.07" />
                    <SPLIT distance="300" swimtime="00:04:02.03" />
                    <SPLIT distance="350" swimtime="00:04:44.13" />
                    <SPLIT distance="400" swimtime="00:05:26.21" />
                    <SPLIT distance="450" swimtime="00:06:07.52" />
                    <SPLIT distance="500" swimtime="00:06:49.31" />
                    <SPLIT distance="550" swimtime="00:07:31.44" />
                    <SPLIT distance="600" swimtime="00:08:13.86" />
                    <SPLIT distance="650" swimtime="00:08:55.35" />
                    <SPLIT distance="700" swimtime="00:09:36.55" />
                    <SPLIT distance="750" swimtime="00:10:16.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="371" swimtime="00:00:29.09" resultid="3838" heatid="10699" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1302" points="389" swimtime="00:01:04.23" resultid="3839" heatid="10779" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="290" swimtime="00:00:33.88" resultid="3840" heatid="10828" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1482" points="345" swimtime="00:02:25.34" resultid="3841" heatid="10860" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:11.35" />
                    <SPLIT distance="150" swimtime="00:01:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="307" swimtime="00:00:39.14" resultid="3842" heatid="10918" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1695" points="345" swimtime="00:05:13.71" resultid="3843" heatid="10941" lane="0" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:15.34" />
                    <SPLIT distance="150" swimtime="00:01:56.59" />
                    <SPLIT distance="200" swimtime="00:02:38.02" />
                    <SPLIT distance="250" swimtime="00:03:18.19" />
                    <SPLIT distance="300" swimtime="00:03:59.11" />
                    <SPLIT distance="350" swimtime="00:04:38.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-24" firstname="Maciej" gender="M" lastname="Brodacki" nation="POL" athleteid="3874">
              <RESULTS>
                <RESULT eventid="1160" points="526" swimtime="00:00:25.90" resultid="3875" heatid="10708" lane="6" entrytime="00:00:26.50" />
                <RESULT eventid="1190" points="432" swimtime="00:02:30.76" resultid="3876" heatid="10729" lane="8" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:09.67" />
                    <SPLIT distance="150" swimtime="00:01:57.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="411" swimtime="00:00:32.33" resultid="3877" heatid="10748" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1302" points="527" swimtime="00:00:58.05" resultid="3878" heatid="10787" lane="7" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="459" swimtime="00:00:29.06" resultid="3879" heatid="10833" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1546" status="DNS" swimtime="00:00:00.00" resultid="3880" heatid="10880" lane="1" entrytime="00:05:45.00" />
                <RESULT eventid="1578" points="425" swimtime="00:01:06.22" resultid="3881" heatid="10891" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="373" swimtime="00:05:05.47" resultid="3882" heatid="10943" lane="7" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:48.67" />
                    <SPLIT distance="200" swimtime="00:02:27.51" />
                    <SPLIT distance="250" swimtime="00:03:06.82" />
                    <SPLIT distance="300" swimtime="00:03:47.53" />
                    <SPLIT distance="350" swimtime="00:04:27.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-07" firstname="Marta" gender="F" lastname="Pachuc" nation="POL" athleteid="3844">
              <RESULTS>
                <RESULT eventid="1144" points="334" swimtime="00:00:34.19" resultid="3845" heatid="10686" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1287" points="325" swimtime="00:01:15.68" resultid="3846" heatid="10770" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="268" swimtime="00:01:39.73" resultid="3847" heatid="10805" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="288" swimtime="00:00:44.63" resultid="3848" heatid="10908" lane="4" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-14" firstname="Kinga" gender="F" lastname="Maciupa" nation="POL" athleteid="3830">
              <RESULTS>
                <RESULT eventid="1175" points="422" swimtime="00:02:48.07" resultid="3831" heatid="10718" lane="1" entrytime="00:02:42.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:18.29" />
                    <SPLIT distance="150" swimtime="00:02:06.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="436" swimtime="00:01:08.61" resultid="3832" heatid="10770" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="408" swimtime="00:00:32.92" resultid="3833" heatid="10823" lane="6" entrytime="00:00:34.32" />
                <RESULT eventid="1437" points="449" swimtime="00:01:15.87" resultid="3834" heatid="10842" lane="5" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="385" swimtime="00:01:16.20" resultid="3835" heatid="10884" lane="3" entrytime="00:01:13.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-20" firstname="Agnieszka" gender="F" lastname="Krzyżostaniak" nation="POL" athleteid="3820">
              <RESULTS>
                <RESULT eventid="1144" points="550" swimtime="00:00:28.95" resultid="3821" heatid="10688" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="1226" points="580" swimtime="00:00:32.44" resultid="3822" heatid="10739" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1287" points="506" swimtime="00:01:05.29" resultid="3823" heatid="10771" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="497" swimtime="00:01:13.33" resultid="3824" heatid="10842" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-09" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="3883">
              <RESULTS>
                <RESULT eventid="1302" points="194" swimtime="00:01:20.98" resultid="3884" heatid="10788" lane="5" entrytime="00:00:54.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-17" firstname="Grzegorz" gender="M" lastname="Juszkiewicz" nation="POL" athleteid="3885">
              <RESULTS>
                <RESULT eventid="1160" points="181" swimtime="00:00:36.96" resultid="3886" heatid="10692" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1242" points="66" swimtime="00:00:59.29" resultid="3887" heatid="10742" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="3888" heatid="10914" lane="1" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-18" firstname="Ola" gender="F" lastname="Szczypek" nation="POL" athleteid="3871">
              <RESULTS>
                <RESULT eventid="1257" points="210" swimtime="00:03:53.84" resultid="3872" heatid="10753" lane="5" entrytime="00:04:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.24" />
                    <SPLIT distance="100" swimtime="00:01:51.68" />
                    <SPLIT distance="150" swimtime="00:02:54.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="206" swimtime="00:01:48.90" resultid="3873" heatid="10805" lane="0" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-19" firstname="Tomasz" gender="M" lastname="Mazur" nation="POL" athleteid="3849">
              <RESULTS>
                <RESULT eventid="1160" points="174" swimtime="00:00:37.44" resultid="3850" heatid="10695" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1302" points="134" swimtime="00:01:31.66" resultid="3851" heatid="10775" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-11-04" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" athleteid="3889">
              <RESULTS>
                <RESULT eventid="1160" points="248" swimtime="00:00:33.26" resultid="3890" heatid="10698" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1242" points="204" swimtime="00:00:40.78" resultid="3891" heatid="10744" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1452" points="179" swimtime="00:01:31.97" resultid="3892" heatid="10846" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="210" swimtime="00:06:10.09" resultid="3893" heatid="10940" lane="9" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                    <SPLIT distance="100" swimtime="00:01:19.62" />
                    <SPLIT distance="150" swimtime="00:02:06.95" />
                    <SPLIT distance="200" swimtime="00:02:54.82" />
                    <SPLIT distance="250" swimtime="00:03:44.28" />
                    <SPLIT distance="300" swimtime="00:04:31.91" />
                    <SPLIT distance="350" swimtime="00:05:22.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-12-12" firstname="Dominika" gender="F" lastname="Zielińska" nation="POL" athleteid="3861">
              <RESULTS>
                <RESULT eventid="1059" points="331" swimtime="00:11:40.59" resultid="3862" heatid="10667" lane="3" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="150" swimtime="00:02:02.65" />
                    <SPLIT distance="200" swimtime="00:02:46.79" />
                    <SPLIT distance="250" swimtime="00:03:31.18" />
                    <SPLIT distance="300" swimtime="00:04:16.76" />
                    <SPLIT distance="350" swimtime="00:05:02.36" />
                    <SPLIT distance="400" swimtime="00:05:47.79" />
                    <SPLIT distance="450" swimtime="00:06:32.42" />
                    <SPLIT distance="500" swimtime="00:07:17.61" />
                    <SPLIT distance="550" swimtime="00:08:02.19" />
                    <SPLIT distance="600" swimtime="00:08:47.66" />
                    <SPLIT distance="650" swimtime="00:09:31.74" />
                    <SPLIT distance="700" swimtime="00:10:16.43" />
                    <SPLIT distance="750" swimtime="00:11:00.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="436" swimtime="00:00:31.29" resultid="3863" heatid="10687" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1175" points="390" swimtime="00:02:52.56" resultid="3864" heatid="10717" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:19.41" />
                    <SPLIT distance="150" swimtime="00:02:09.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="368" swimtime="00:00:37.75" resultid="3865" heatid="10738" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1287" points="427" swimtime="00:01:09.12" resultid="3866" heatid="10770" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat C  35-39  lat" eventid="1437" points="409" swimtime="00:01:18.26" resultid="3867" heatid="10841" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="381" swimtime="00:02:35.73" resultid="3868" heatid="10855" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:16.87" />
                    <SPLIT distance="150" swimtime="00:01:57.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="339" swimtime="00:01:19.52" resultid="3869" heatid="10884" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1593" points="397" swimtime="00:02:48.76" resultid="3870" heatid="10897" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                    <SPLIT distance="100" swimtime="00:01:22.71" />
                    <SPLIT distance="150" swimtime="00:02:06.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="348" swimtime="00:02:12.79" resultid="3897" heatid="10801" lane="1" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:09.22" />
                    <SPLIT distance="150" swimtime="00:01:43.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3874" number="1" />
                    <RELAYPOSITION athleteid="3825" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3852" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3836" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" points="419" swimtime="00:01:53.33" resultid="3898" heatid="10872" lane="9" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:00:59.24" />
                    <SPLIT distance="150" swimtime="00:01:27.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3852" number="1" />
                    <RELAYPOSITION athleteid="3836" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3825" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3874" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1518" points="212" status="EXH" swimtime="00:02:22.20" resultid="3901" heatid="10870" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:49.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3883" number="1" />
                    <RELAYPOSITION athleteid="3885" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3849" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3889" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1347" points="399" status="EXH" swimtime="00:02:24.34" resultid="3899" heatid="10798" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="150" swimtime="00:01:53.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3820" number="1" />
                    <RELAYPOSITION athleteid="3871" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3830" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3861" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1497" points="343" status="EXH" swimtime="00:02:17.89" resultid="3900" heatid="10868" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="100" swimtime="00:01:14.40" />
                    <SPLIT distance="150" swimtime="00:01:46.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3861" number="1" />
                    <RELAYPOSITION athleteid="3871" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3844" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3830" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:01:58.88" resultid="3894" heatid="10733" lane="3" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.95" />
                    <SPLIT distance="100" swimtime="00:00:59.05" />
                    <SPLIT distance="150" swimtime="00:01:32.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3825" number="1" />
                    <RELAYPOSITION athleteid="3861" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3844" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3874" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1653" swimtime="00:02:16.18" resultid="3895" heatid="10929" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                    <SPLIT distance="150" swimtime="00:01:50.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3844" number="1" />
                    <RELAYPOSITION athleteid="3825" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3861" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3874" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1205" status="EXH" swimtime="00:02:04.83" resultid="3896" heatid="10733" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:02.99" />
                    <SPLIT distance="150" swimtime="00:01:35.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3852" number="1" />
                    <RELAYPOSITION athleteid="3830" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3889" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3820" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SWPRA" nation="CZE" clubid="2938" name="Swimmpower Prague">
          <CONTACT city="Prague" email="info@swim.by" name="Swimmpower Prague, z.s." phone="+375291555114" street="Luzicka 9" />
          <ATHLETES>
            <ATHLETE birthdate="1983-05-01" firstname="Andrzej" gender="M" lastname="Waszkewicz" nation="POL" athleteid="2946">
              <RESULTS>
                <RESULT eventid="1160" points="590" swimtime="00:00:24.92" resultid="7908" heatid="10711" lane="2" entrytime="00:00:24.41" entrycourse="LCM" />
                <RESULT eventid="1422" points="609" swimtime="00:00:26.46" resultid="7909" heatid="10838" lane="1" entrytime="00:00:26.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Andrea" gender="F" lastname="Janigova" nation="CZE" athleteid="9532">
              <RESULTS>
                <RESULT eventid="1257" points="330" swimtime="00:03:21.25" resultid="9533" heatid="10756" lane="0" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                    <SPLIT distance="100" swimtime="00:01:38.04" />
                    <SPLIT distance="150" swimtime="00:02:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="332" swimtime="00:01:32.84" resultid="9534" heatid="10808" lane="0" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="347" swimtime="00:00:41.92" resultid="9535" heatid="10910" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAOPO" nation="POL" region="OPO" clubid="4513" name="T.P.Masters Opole">
          <CONTACT city="OPOLE" email="OPOLBUD@ONET.EU" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Witkowski" nation="POL" athleteid="4540">
              <RESULTS>
                <RESULT eventid="1160" points="107" swimtime="00:00:44.04" resultid="7749" heatid="10692" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1242" points="73" swimtime="00:00:57.43" resultid="7750" heatid="10741" lane="3" entrytime="00:00:56.00" />
                <RESULT eventid="1302" points="61" swimtime="00:01:58.67" resultid="7751" heatid="10774" lane="9" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="40" swimtime="00:02:30.55" resultid="7752" heatid="10844" lane="7" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="7753" heatid="10857" lane="8" entrytime="00:03:59.00" />
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="7754" heatid="10899" lane="4" entrytime="00:04:35.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="7755" heatid="10913" lane="2" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Tomasz" gender="M" lastname="Samsel" nation="POL" athleteid="4527">
              <RESULTS>
                <RESULT eventid="1098" points="323" swimtime="00:10:58.56" resultid="7738" heatid="10672" lane="7" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:50.88" />
                    <SPLIT distance="200" swimtime="00:02:31.06" />
                    <SPLIT distance="250" swimtime="00:03:11.87" />
                    <SPLIT distance="300" swimtime="00:03:52.76" />
                    <SPLIT distance="350" swimtime="00:04:34.35" />
                    <SPLIT distance="400" swimtime="00:05:16.84" />
                    <SPLIT distance="450" swimtime="00:05:59.65" />
                    <SPLIT distance="500" swimtime="00:06:42.52" />
                    <SPLIT distance="550" swimtime="00:07:26.02" />
                    <SPLIT distance="600" swimtime="00:08:09.77" />
                    <SPLIT distance="650" swimtime="00:08:53.64" />
                    <SPLIT distance="700" swimtime="00:09:36.63" />
                    <SPLIT distance="750" swimtime="00:10:19.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="492" swimtime="00:00:26.47" resultid="7739" heatid="10709" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1302" points="517" swimtime="00:00:58.44" resultid="7740" heatid="10787" lane="8" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="334" swimtime="00:00:32.32" resultid="7741" heatid="10834" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1482" points="426" swimtime="00:02:15.51" resultid="7742" heatid="10865" lane="8" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:07.28" />
                    <SPLIT distance="150" swimtime="00:01:42.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="7743" heatid="10888" lane="3" entrytime="00:01:16.00" />
                <RESULT eventid="1695" points="369" swimtime="00:05:06.68" resultid="7744" heatid="10943" lane="1" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:13.13" />
                    <SPLIT distance="150" swimtime="00:01:53.39" />
                    <SPLIT distance="200" swimtime="00:02:33.84" />
                    <SPLIT distance="250" swimtime="00:03:13.32" />
                    <SPLIT distance="300" swimtime="00:03:52.24" />
                    <SPLIT distance="350" swimtime="00:04:30.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Zbigniew" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="4535">
              <RESULTS>
                <RESULT eventid="1190" points="403" swimtime="00:02:34.25" resultid="7745" heatid="10727" lane="3" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:09.83" />
                    <SPLIT distance="150" swimtime="00:01:58.43" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn  w  kat G  55-59  lat" eventid="1242" points="426" swimtime="00:00:31.94" resultid="7746" heatid="10749" lane="4" entrytime="00:00:31.20" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn w  kat G 55-59  lat" eventid="1452" points="437" swimtime="00:01:08.29" resultid="7747" heatid="10850" lane="9" entrytime="00:01:06.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1608" points="433" swimtime="00:02:27.93" resultid="7748" heatid="10904" lane="2" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:01:50.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Bartnikowska" nation="POL" athleteid="4548">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat A 25-29 lat" eventid="1113" points="350" swimtime="00:21:52.04" resultid="7756" heatid="10674" lane="3" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:20.63" />
                    <SPLIT distance="150" swimtime="00:02:04.01" />
                    <SPLIT distance="200" swimtime="00:02:47.94" />
                    <SPLIT distance="250" swimtime="00:03:32.85" />
                    <SPLIT distance="300" swimtime="00:04:17.20" />
                    <SPLIT distance="350" swimtime="00:05:01.43" />
                    <SPLIT distance="400" swimtime="00:05:45.38" />
                    <SPLIT distance="450" swimtime="00:06:29.83" />
                    <SPLIT distance="500" swimtime="00:07:13.75" />
                    <SPLIT distance="550" swimtime="00:07:58.42" />
                    <SPLIT distance="600" swimtime="00:08:43.19" />
                    <SPLIT distance="650" swimtime="00:09:27.86" />
                    <SPLIT distance="700" swimtime="00:10:11.93" />
                    <SPLIT distance="750" swimtime="00:10:56.42" />
                    <SPLIT distance="800" swimtime="00:11:40.19" />
                    <SPLIT distance="850" swimtime="00:12:24.80" />
                    <SPLIT distance="900" swimtime="00:13:09.34" />
                    <SPLIT distance="950" swimtime="00:13:53.83" />
                    <SPLIT distance="1000" swimtime="00:14:37.94" />
                    <SPLIT distance="1050" swimtime="00:15:22.29" />
                    <SPLIT distance="1100" swimtime="00:16:06.15" />
                    <SPLIT distance="1150" swimtime="00:16:50.70" />
                    <SPLIT distance="1200" swimtime="00:17:34.84" />
                    <SPLIT distance="1250" swimtime="00:18:15.77" />
                    <SPLIT distance="1300" swimtime="00:19:03.81" />
                    <SPLIT distance="1350" swimtime="00:19:48.29" />
                    <SPLIT distance="1400" swimtime="00:20:31.54" />
                    <SPLIT distance="1450" swimtime="00:21:13.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="484" swimtime="00:00:30.22" resultid="7757" heatid="10687" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1175" points="472" swimtime="00:02:41.94" resultid="7758" heatid="10717" lane="2" entrytime="00:02:49.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="100" swimtime="00:01:17.18" />
                    <SPLIT distance="150" swimtime="00:02:05.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="521" swimtime="00:00:33.62" resultid="7759" heatid="10738" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1407" points="460" swimtime="00:00:31.63" resultid="7760" heatid="10824" lane="9" entrytime="00:00:33.53" />
                <RESULT eventid="1525" points="419" swimtime="00:05:55.92" resultid="7761" heatid="10875" lane="0" entrytime="00:06:06.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                    <SPLIT distance="100" swimtime="00:01:28.10" />
                    <SPLIT distance="150" swimtime="00:02:11.82" />
                    <SPLIT distance="200" swimtime="00:02:55.77" />
                    <SPLIT distance="250" swimtime="00:03:49.03" />
                    <SPLIT distance="300" swimtime="00:04:39.08" />
                    <SPLIT distance="350" swimtime="00:05:19.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="463" swimtime="00:02:40.30" resultid="7762" heatid="10897" lane="6" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:20.35" />
                    <SPLIT distance="150" swimtime="00:02:01.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AQBAR" nation="POL" region="WIE" clubid="3794" name="Team Masters Aquapark Barracuda" shortname="Team Masters Aquapark Barracud">
          <CONTACT city="KALISZ" email="galczynskiwoj@op.pl" name="GAŁCZYŃSKI WOJCIECH" phone="790690666" state="WLKP" street="PODMIEJSKA 15/28" zip="62-800" />
          <ATHLETES>
            <ATHLETE birthdate="1986-07-20" firstname="Mateusz" gender="M" lastname="Szuleta" nation="POL" athleteid="3802">
              <RESULTS>
                <RESULT eventid="1160" points="381" swimtime="00:00:28.82" resultid="6302" heatid="10708" lane="9" entrytime="00:00:27.00" />
                <RESULT eventid="1392" points="327" swimtime="00:01:22.85" resultid="6303" heatid="10818" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="436" swimtime="00:00:34.83" resultid="6304" heatid="10925" lane="7" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-09-12" firstname="Wojciech" gender="M" lastname="Gałczyński" nation="POL" athleteid="3795">
              <RESULTS>
                <RESULT eventid="1160" points="487" swimtime="00:00:26.56" resultid="6296" heatid="10707" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1242" points="372" swimtime="00:00:33.40" resultid="6297" heatid="10748" lane="6" entrytime="00:00:33.55" />
                <RESULT eventid="1272" points="343" swimtime="00:03:01.27" resultid="6298" heatid="10762" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:23.53" />
                    <SPLIT distance="150" swimtime="00:02:10.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="394" swimtime="00:01:17.89" resultid="6299" heatid="10818" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="321" swimtime="00:01:15.65" resultid="6300" heatid="10848" lane="0" entrytime="00:01:16.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="487" swimtime="00:00:33.56" resultid="6301" heatid="10925" lane="9" entrytime="00:00:33.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-01" firstname="Andrzej" gender="M" lastname="Sypniewski" nation="POL" athleteid="3806">
              <RESULTS>
                <RESULT eventid="1190" points="218" swimtime="00:03:09.28" resultid="6305" heatid="10722" lane="1" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                    <SPLIT distance="100" swimtime="00:01:28.53" />
                    <SPLIT distance="150" swimtime="00:02:21.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="229" swimtime="00:03:27.56" resultid="6306" heatid="10760" lane="5" entrytime="00:03:18.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.59" />
                    <SPLIT distance="100" swimtime="00:01:39.53" />
                    <SPLIT distance="150" swimtime="00:02:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="125" swimtime="00:03:43.00" resultid="6307" heatid="10792" lane="4" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:39.64" />
                    <SPLIT distance="150" swimtime="00:02:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="229" swimtime="00:01:33.27" resultid="6308" heatid="10813" lane="4" entrytime="00:01:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="181" swimtime="00:07:10.51" resultid="6309" heatid="10878" lane="9" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.04" />
                    <SPLIT distance="100" swimtime="00:01:41.87" />
                    <SPLIT distance="150" swimtime="00:02:37.74" />
                    <SPLIT distance="200" swimtime="00:03:33.07" />
                    <SPLIT distance="250" swimtime="00:04:31.00" />
                    <SPLIT distance="300" swimtime="00:05:30.83" />
                    <SPLIT distance="350" swimtime="00:06:21.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="128" swimtime="00:01:38.75" resultid="6310" heatid="10886" lane="4" entrytime="00:01:32.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="262" swimtime="00:00:41.27" resultid="6311" heatid="10917" lane="5" entrytime="00:00:40.21" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5130" nation="GER" region="17" clubid="3472" name="TG Lage 1862">
          <CONTACT city="Lage" email="tg-schwimmen@gmx.de" name="Ute Lange" state="NO" street="Ringstrasse 3" zip="32791" />
          <ATHLETES>
            <ATHLETE birthdate="1968-04-07" firstname="Konstantin" gender="M" lastname="Sklyar" nation="GER" license="321129" athleteid="3473">
              <RESULTS>
                <RESULT eventid="1098" points="328" swimtime="00:10:55.05" resultid="8296" heatid="10671" lane="1" entrytime="00:11:31.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:56.58" />
                    <SPLIT distance="200" swimtime="00:02:38.24" />
                    <SPLIT distance="250" swimtime="00:03:19.59" />
                    <SPLIT distance="300" swimtime="00:04:01.52" />
                    <SPLIT distance="350" swimtime="00:04:43.14" />
                    <SPLIT distance="400" swimtime="00:05:25.19" />
                    <SPLIT distance="450" swimtime="00:06:06.66" />
                    <SPLIT distance="500" swimtime="00:06:48.71" />
                    <SPLIT distance="550" swimtime="00:07:30.22" />
                    <SPLIT distance="600" swimtime="00:08:12.10" />
                    <SPLIT distance="650" swimtime="00:08:53.29" />
                    <SPLIT distance="700" swimtime="00:09:35.10" />
                    <SPLIT distance="750" swimtime="00:10:15.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="8297" heatid="10761" lane="2" entrytime="00:03:09.88" entrycourse="LCM" />
                <RESULT eventid="1332" status="DNS" swimtime="00:00:00.00" resultid="8298" heatid="10794" lane="1" entrytime="00:03:01.50" entrycourse="LCM" />
                <RESULT eventid="1482" points="309" swimtime="00:02:30.81" resultid="8299" heatid="10861" lane="5" entrytime="00:02:28.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:51.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="273" swimtime="00:06:15.85" resultid="8300" heatid="10879" lane="6" entrytime="00:06:08.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                    <SPLIT distance="100" swimtime="00:01:24.74" />
                    <SPLIT distance="150" swimtime="00:02:14.54" />
                    <SPLIT distance="200" swimtime="00:03:03.57" />
                    <SPLIT distance="250" swimtime="00:03:58.08" />
                    <SPLIT distance="300" swimtime="00:04:52.64" />
                    <SPLIT distance="350" swimtime="00:05:34.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="8301" heatid="10889" lane="8" entrytime="00:01:14.11" entrycourse="LCM" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="8302" heatid="10942" lane="2" entrytime="00:05:11.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ALVSE" nation="CZE" clubid="3058" name="TJ Alcedo Vsetín z.s.">
          <CONTACT city="Vsetín" email="pavel.obr@czechswimming.cz" name="Pavel Obr" phone="+420724955185" state="CZE" street="Dolní Jasenka 770" zip="755 01" />
          <ATHLETES>
            <ATHLETE birthdate="1967-05-03" firstname="Pavel" gender="M" lastname="Obr" nation="CZE" athleteid="3087">
              <RESULTS>
                <RESULT eventid="1160" points="424" swimtime="00:00:27.82" resultid="6282" heatid="10704" lane="4" entrytime="00:00:28.16" />
                <RESULT eventid="1190" points="343" swimtime="00:02:42.83" resultid="6283" heatid="10726" lane="5" entrytime="00:02:40.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:15.14" />
                    <SPLIT distance="150" swimtime="00:02:03.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="434" swimtime="00:01:01.94" resultid="6284" heatid="10783" lane="5" entrytime="00:01:02.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="440" swimtime="00:00:29.47" resultid="6285" heatid="10833" lane="3" entrytime="00:00:30.76" />
                <RESULT eventid="1546" points="280" swimtime="00:06:12.39" resultid="6286" heatid="10879" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:19.36" />
                    <SPLIT distance="150" swimtime="00:02:09.96" />
                    <SPLIT distance="200" swimtime="00:03:00.58" />
                    <SPLIT distance="250" swimtime="00:03:52.27" />
                    <SPLIT distance="300" swimtime="00:04:46.14" />
                    <SPLIT distance="350" swimtime="00:05:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="390" swimtime="00:00:36.16" resultid="6287" heatid="10921" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-04-15" firstname="Bronislava" gender="F" lastname="Kudelová" nation="CZE" athleteid="3094">
              <RESULTS>
                <RESULT eventid="1175" points="251" swimtime="00:03:19.93" resultid="6288" heatid="10716" lane="0" entrytime="00:03:09.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:01:33.87" />
                    <SPLIT distance="150" swimtime="00:02:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="296" swimtime="00:00:40.58" resultid="6289" heatid="10737" lane="4" entrytime="00:00:38.90" />
                <RESULT eventid="1437" points="264" swimtime="00:01:30.54" resultid="6291" heatid="10841" lane="1" entrytime="00:01:28.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="229" swimtime="00:07:15.19" resultid="6292" heatid="10874" lane="1" entrytime="00:06:57.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                    <SPLIT distance="100" swimtime="00:01:41.25" />
                    <SPLIT distance="150" swimtime="00:02:36.47" />
                    <SPLIT distance="200" swimtime="00:03:30.85" />
                    <SPLIT distance="250" swimtime="00:04:31.75" />
                    <SPLIT distance="300" swimtime="00:05:34.33" />
                    <SPLIT distance="350" swimtime="00:06:25.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="250" swimtime="00:03:16.80" resultid="6293" heatid="10896" lane="7" entrytime="00:03:08.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                    <SPLIT distance="100" swimtime="00:01:34.51" />
                    <SPLIT distance="150" swimtime="00:02:26.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="311" swimtime="00:00:35.00" resultid="10652" heatid="10680" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKOS" nation="POL" region="ZAC" clubid="4914" name="Tkkf Koszalin Masters">
          <CONTACT city="Koszalin" email="jakubkielar3@gmail.com" name="Kielar" />
          <ATHLETES>
            <ATHLETE birthdate="1974-06-28" firstname="Michał" gender="M" lastname="Pieślak" nation="POL" athleteid="4921">
              <RESULTS>
                <RESULT eventid="1160" points="406" swimtime="00:00:28.23" resultid="6576" heatid="10702" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1302" points="374" swimtime="00:01:05.10" resultid="6577" heatid="10781" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="280" swimtime="00:01:27.24" resultid="6578" heatid="10814" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="325" swimtime="00:02:28.24" resultid="6579" heatid="10862" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:09.37" />
                    <SPLIT distance="150" swimtime="00:01:47.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="334" swimtime="00:00:38.07" resultid="6580" heatid="10919" lane="4" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-05" firstname="Agnieszka" gender="F" lastname="Paziewska" nation="POL" athleteid="4927">
              <RESULTS>
                <RESULT eventid="1144" points="341" swimtime="00:00:33.95" resultid="6581" heatid="10686" lane="1" entrytime="00:00:33.50" />
                <RESULT eventid="1287" points="308" swimtime="00:01:17.05" resultid="6582" heatid="10769" lane="9" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="6583" heatid="10805" lane="5" entrytime="00:01:41.00" />
                <RESULT eventid="1467" points="284" swimtime="00:02:51.83" resultid="6584" heatid="10853" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:23.56" />
                    <SPLIT distance="150" swimtime="00:02:09.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="262" swimtime="00:00:46.05" resultid="6585" heatid="10909" lane="8" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-22" firstname="Grzegorz" gender="M" lastname="Ćwikła" nation="POL" athleteid="4915">
              <RESULTS>
                <RESULT eventid="1128" points="279" swimtime="00:22:12.21" resultid="6571" heatid="10677" lane="3" entrytime="00:22:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:19.31" />
                    <SPLIT distance="150" swimtime="00:02:02.79" />
                    <SPLIT distance="200" swimtime="00:02:46.84" />
                    <SPLIT distance="250" swimtime="00:03:30.95" />
                    <SPLIT distance="300" swimtime="00:04:15.02" />
                    <SPLIT distance="350" swimtime="00:04:59.33" />
                    <SPLIT distance="400" swimtime="00:05:43.59" />
                    <SPLIT distance="450" swimtime="00:06:27.95" />
                    <SPLIT distance="500" swimtime="00:07:12.70" />
                    <SPLIT distance="550" swimtime="00:07:57.46" />
                    <SPLIT distance="600" swimtime="00:08:42.44" />
                    <SPLIT distance="650" swimtime="00:09:27.00" />
                    <SPLIT distance="700" swimtime="00:10:12.13" />
                    <SPLIT distance="750" swimtime="00:10:57.54" />
                    <SPLIT distance="800" swimtime="00:11:42.97" />
                    <SPLIT distance="850" swimtime="00:12:28.73" />
                    <SPLIT distance="900" swimtime="00:13:14.24" />
                    <SPLIT distance="950" swimtime="00:14:00.06" />
                    <SPLIT distance="1000" swimtime="00:14:45.51" />
                    <SPLIT distance="1050" swimtime="00:15:30.82" />
                    <SPLIT distance="1100" swimtime="00:16:16.20" />
                    <SPLIT distance="1150" swimtime="00:17:01.55" />
                    <SPLIT distance="1200" swimtime="00:17:47.43" />
                    <SPLIT distance="1250" swimtime="00:18:33.02" />
                    <SPLIT distance="1300" swimtime="00:19:18.71" />
                    <SPLIT distance="1350" swimtime="00:20:04.10" />
                    <SPLIT distance="1400" swimtime="00:20:49.43" />
                    <SPLIT distance="1450" swimtime="00:21:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="288" swimtime="00:01:18.50" resultid="6572" heatid="10848" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="277" swimtime="00:06:13.83" resultid="6573" heatid="10879" lane="0" entrytime="00:06:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:25.24" />
                    <SPLIT distance="150" swimtime="00:02:17.80" />
                    <SPLIT distance="200" swimtime="00:03:07.59" />
                    <SPLIT distance="250" swimtime="00:04:03.35" />
                    <SPLIT distance="300" swimtime="00:04:57.16" />
                    <SPLIT distance="350" swimtime="00:05:36.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="266" swimtime="00:02:54.01" resultid="6574" heatid="10902" lane="3" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:26.62" />
                    <SPLIT distance="150" swimtime="00:02:11.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="299" swimtime="00:05:28.76" resultid="6575" heatid="10942" lane="0" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="100" swimtime="00:01:16.90" />
                    <SPLIT distance="150" swimtime="00:01:58.82" />
                    <SPLIT distance="200" swimtime="00:02:41.83" />
                    <SPLIT distance="250" swimtime="00:03:25.01" />
                    <SPLIT distance="300" swimtime="00:04:08.57" />
                    <SPLIT distance="350" swimtime="00:04:50.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-29" firstname="Lidia" gender="F" lastname="Mikołajczyk" nation="POL" athleteid="4938">
              <RESULTS>
                <RESULT eventid="1175" points="346" swimtime="00:02:59.58" resultid="6590" heatid="10717" lane="9" entrytime="00:02:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:23.24" />
                    <SPLIT distance="150" swimtime="00:02:15.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="314" swimtime="00:03:24.58" resultid="6591" heatid="10755" lane="3" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:36.98" />
                    <SPLIT distance="150" swimtime="00:02:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="336" swimtime="00:01:32.55" resultid="6592" heatid="10807" lane="8" entrytime="00:01:31.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="307" swimtime="00:06:34.47" resultid="6593" heatid="10874" lane="4" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="100" swimtime="00:01:32.56" />
                    <SPLIT distance="150" swimtime="00:02:23.71" />
                    <SPLIT distance="200" swimtime="00:03:13.87" />
                    <SPLIT distance="250" swimtime="00:04:07.99" />
                    <SPLIT distance="300" swimtime="00:05:04.04" />
                    <SPLIT distance="350" swimtime="00:05:50.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="6594" heatid="10910" lane="0" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-24" firstname="Wioletta" gender="F" lastname="Pawliczek" nation="POL" athleteid="4933">
              <RESULTS>
                <RESULT eventid="1144" points="284" swimtime="00:00:36.08" resultid="6586" heatid="10684" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1226" points="310" swimtime="00:00:39.96" resultid="6587" heatid="10736" lane="6" entrytime="00:00:43.61" />
                <RESULT eventid="1437" points="284" swimtime="00:01:28.37" resultid="6588" heatid="10841" lane="8" entrytime="00:01:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="255" swimtime="00:03:15.58" resultid="6589" heatid="10895" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.73" />
                    <SPLIT distance="100" swimtime="00:01:37.06" />
                    <SPLIT distance="150" swimtime="00:02:28.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:23.60" resultid="6595" heatid="10927" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.23" />
                    <SPLIT distance="150" swimtime="00:01:54.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4933" number="1" />
                    <RELAYPOSITION athleteid="4938" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4915" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4921" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TORPE" nation="LTU" clubid="3481" name="Torpedos">
          <CONTACT email="vilmantasenator@gmail.com" name="Vilmantas Krasauskas" phone="+37068746068" />
          <ATHLETES>
            <ATHLETE birthdate="1964-07-31" firstname="Vilmantas" gender="M" lastname="Krasauskas" nation="LTU" athleteid="3501">
              <RESULTS>
                <RESULT eventid="1302" points="379" swimtime="00:01:04.80" resultid="8320" heatid="10783" lane="8" entrytime="00:01:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="354" swimtime="00:02:24.12" resultid="8321" heatid="10862" lane="5" entrytime="00:02:22.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:46.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="8322" heatid="10942" lane="4" entrytime="00:05:07.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-04" firstname="Jurate" gender="F" lastname="Pranckeviciene" nation="LTU" athleteid="3482">
              <RESULTS>
                <RESULT eventid="1226" status="DNS" swimtime="00:00:00.00" resultid="8304" heatid="10736" lane="0" entrytime="00:00:46.00" entrycourse="LCM" />
                <RESULT eventid="1287" points="310" swimtime="00:01:16.92" resultid="8305" heatid="10769" lane="1" entrytime="00:01:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="227" swimtime="00:00:40.00" resultid="8306" heatid="10821" lane="4" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1467" points="237" swimtime="00:03:02.43" resultid="8307" heatid="10853" lane="1" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:01:28.92" />
                    <SPLIT distance="150" swimtime="00:02:17.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="192" swimtime="00:03:34.72" resultid="8308" heatid="10895" lane="3" entrytime="00:03:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.85" />
                    <SPLIT distance="100" swimtime="00:01:44.36" />
                    <SPLIT distance="150" swimtime="00:02:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" status="DNS" swimtime="00:00:00.00" resultid="8309" heatid="10933" lane="9" entrytime="00:06:20.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-02-07" firstname="Margarita" gender="F" lastname="Cineliene" nation="LTU" athleteid="3489">
              <RESULTS>
                <RESULT eventid="1257" points="188" swimtime="00:04:02.54" resultid="8310" heatid="10754" lane="6" entrytime="00:03:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                    <SPLIT distance="100" swimtime="00:01:56.28" />
                    <SPLIT distance="150" swimtime="00:02:59.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="204" swimtime="00:01:49.17" resultid="8311" heatid="10805" lane="9" entrytime="00:01:48.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="93" swimtime="00:00:53.83" resultid="8312" heatid="10821" lane="9" entrytime="00:00:54.00" entrycourse="LCM" />
                <RESULT eventid="1623" points="235" swimtime="00:00:47.76" resultid="8313" heatid="10907" lane="4" entrytime="00:00:48.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-03-14" firstname="Stasys" gender="M" lastname="Grigas" nation="LTU" athleteid="3494">
              <RESULTS>
                <RESULT eventid="1242" points="53" swimtime="00:01:03.88" resultid="8314" heatid="10744" lane="9" entrytime="00:01:03.00" entrycourse="LCM" />
                <RESULT eventid="1302" points="46" swimtime="00:02:10.70" resultid="8315" heatid="10773" lane="2" entrytime="00:02:09.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="48" swimtime="00:02:21.74" resultid="8316" heatid="10844" lane="8" entrytime="00:02:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="31" swimtime="00:05:21.90" resultid="8317" heatid="10856" lane="4" entrytime="00:05:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.53" />
                    <SPLIT distance="100" swimtime="00:02:42.37" />
                    <SPLIT distance="150" swimtime="00:04:03.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="47" swimtime="00:05:09.81" resultid="8318" heatid="10899" lane="2" entrytime="00:05:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.76" />
                    <SPLIT distance="100" swimtime="00:02:34.65" />
                    <SPLIT distance="150" swimtime="00:03:55.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="92" swimtime="00:00:58.41" resultid="8319" heatid="10913" lane="6" entrytime="00:00:59.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02602" nation="POL" region="KUJ" clubid="3902" name="Toruń Multisport Team">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="3924">
              <RESULTS>
                <RESULT eventid="1098" points="185" swimtime="00:13:12.49" resultid="8331" heatid="10670" lane="2" entrytime="00:12:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.50" />
                    <SPLIT distance="100" swimtime="00:01:35.16" />
                    <SPLIT distance="150" swimtime="00:02:25.28" />
                    <SPLIT distance="200" swimtime="00:03:17.29" />
                    <SPLIT distance="250" swimtime="00:04:07.95" />
                    <SPLIT distance="300" swimtime="00:04:59.29" />
                    <SPLIT distance="350" swimtime="00:05:50.17" />
                    <SPLIT distance="400" swimtime="00:06:40.52" />
                    <SPLIT distance="450" swimtime="00:07:31.87" />
                    <SPLIT distance="500" swimtime="00:08:22.77" />
                    <SPLIT distance="550" swimtime="00:09:12.77" />
                    <SPLIT distance="600" swimtime="00:10:03.76" />
                    <SPLIT distance="650" swimtime="00:10:53.24" />
                    <SPLIT distance="700" swimtime="00:11:43.93" />
                    <SPLIT distance="750" swimtime="00:12:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="264" swimtime="00:00:32.56" resultid="8332" heatid="10697" lane="4" entrytime="00:00:32.30" />
                <RESULT eventid="1302" points="249" swimtime="00:01:14.50" resultid="8333" heatid="10778" lane="2" entrytime="00:01:11.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="219" swimtime="00:00:37.20" resultid="8334" heatid="10829" lane="0" entrytime="00:00:36.50" />
                <RESULT eventid="1482" points="200" swimtime="00:02:54.35" resultid="8335" heatid="10860" lane="8" entrytime="00:02:48.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:01:26.65" />
                    <SPLIT distance="150" swimtime="00:02:13.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="142" swimtime="00:01:35.47" resultid="8336" heatid="10887" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-08-21" firstname="Tomasz" gender="M" lastname="Osóbka" nation="POL" athleteid="3946">
              <RESULTS>
                <RESULT eventid="1160" points="35" swimtime="00:01:03.82" resultid="8350" heatid="10690" lane="5" entrytime="00:01:04.56" />
                <RESULT eventid="1302" points="13" swimtime="00:03:18.48" resultid="8351" heatid="10773" lane="1" entrytime="00:02:31.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="8352" heatid="10809" lane="6" entrytime="00:02:58.00" />
                <RESULT eventid="1638" points="22" swimtime="00:01:34.25" resultid="8353" heatid="10912" lane="4" entrytime="00:01:28.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-10-23" firstname="Marcin" gender="M" lastname="Mykowski" nation="POL" athleteid="3919">
              <RESULTS>
                <RESULT eventid="1098" points="329" swimtime="00:10:54.41" resultid="8327" heatid="10671" lane="9" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:14.93" />
                    <SPLIT distance="150" swimtime="00:01:56.13" />
                    <SPLIT distance="200" swimtime="00:02:37.67" />
                    <SPLIT distance="250" swimtime="00:03:20.61" />
                    <SPLIT distance="300" swimtime="00:04:03.03" />
                    <SPLIT distance="350" swimtime="00:04:45.91" />
                    <SPLIT distance="400" swimtime="00:05:28.15" />
                    <SPLIT distance="450" swimtime="00:06:09.87" />
                    <SPLIT distance="500" swimtime="00:06:52.00" />
                    <SPLIT distance="550" swimtime="00:07:34.03" />
                    <SPLIT distance="600" swimtime="00:08:16.43" />
                    <SPLIT distance="650" swimtime="00:08:56.68" />
                    <SPLIT distance="700" swimtime="00:09:36.93" />
                    <SPLIT distance="750" swimtime="00:10:16.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="484" swimtime="00:00:59.74" resultid="8328" heatid="10781" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="362" swimtime="00:02:23.05" resultid="8329" heatid="10863" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:10.00" />
                    <SPLIT distance="150" swimtime="00:01:47.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="8330" heatid="10902" lane="2" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="3951">
              <RESULTS>
                <RESULT eventid="1190" points="51" swimtime="00:05:07.26" resultid="8354" heatid="10719" lane="6" entrytime="00:05:01.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.89" />
                    <SPLIT distance="100" swimtime="00:02:37.92" />
                    <SPLIT distance="150" swimtime="00:04:10.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="39" swimtime="00:01:10.41" resultid="8355" heatid="10741" lane="9" entrytime="00:01:10.83" />
                <RESULT eventid="1332" status="DNS" swimtime="00:00:00.00" resultid="8356" heatid="10791" lane="3" entrytime="00:05:46.80" />
                <RESULT eventid="1482" points="73" swimtime="00:04:03.44" resultid="8357" heatid="10857" lane="9" entrytime="00:04:00.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.42" />
                    <SPLIT distance="100" swimtime="00:01:58.97" />
                    <SPLIT distance="150" swimtime="00:03:00.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="50" swimtime="00:10:59.97" resultid="8358" heatid="10876" lane="6" entrytime="00:10:38.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.01" />
                    <SPLIT distance="100" swimtime="00:02:44.02" />
                    <SPLIT distance="150" swimtime="00:04:21.63" />
                    <SPLIT distance="200" swimtime="00:05:42.26" />
                    <SPLIT distance="250" swimtime="00:07:21.85" />
                    <SPLIT distance="300" swimtime="00:08:56.43" />
                    <SPLIT distance="350" swimtime="00:09:59.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="32" swimtime="00:02:35.34" resultid="8359" heatid="10885" lane="2" entrytime="00:02:34.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="33" swimtime="00:05:47.15" resultid="8360" heatid="10899" lane="6" entrytime="00:05:28.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.90" />
                    <SPLIT distance="100" swimtime="00:02:55.36" />
                    <SPLIT distance="150" swimtime="00:04:23.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-28" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="3967">
              <RESULTS>
                <RESULT eventid="1128" points="399" swimtime="00:19:42.63" resultid="8368" heatid="10679" lane="3" entrytime="00:19:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:47.33" />
                    <SPLIT distance="200" swimtime="00:02:25.90" />
                    <SPLIT distance="250" swimtime="00:03:04.83" />
                    <SPLIT distance="300" swimtime="00:03:44.49" />
                    <SPLIT distance="350" swimtime="00:04:24.17" />
                    <SPLIT distance="400" swimtime="00:05:04.38" />
                    <SPLIT distance="450" swimtime="00:05:44.40" />
                    <SPLIT distance="500" swimtime="00:06:24.77" />
                    <SPLIT distance="550" swimtime="00:07:05.06" />
                    <SPLIT distance="600" swimtime="00:07:45.29" />
                    <SPLIT distance="650" swimtime="00:08:25.86" />
                    <SPLIT distance="700" swimtime="00:09:06.46" />
                    <SPLIT distance="750" swimtime="00:09:46.64" />
                    <SPLIT distance="800" swimtime="00:10:26.79" />
                    <SPLIT distance="850" swimtime="00:11:06.80" />
                    <SPLIT distance="900" swimtime="00:11:47.12" />
                    <SPLIT distance="950" swimtime="00:12:27.34" />
                    <SPLIT distance="1000" swimtime="00:13:07.50" />
                    <SPLIT distance="1050" swimtime="00:13:47.83" />
                    <SPLIT distance="1100" swimtime="00:14:28.10" />
                    <SPLIT distance="1150" swimtime="00:15:08.44" />
                    <SPLIT distance="1200" swimtime="00:15:48.61" />
                    <SPLIT distance="1250" swimtime="00:16:28.95" />
                    <SPLIT distance="1300" swimtime="00:17:08.77" />
                    <SPLIT distance="1350" swimtime="00:17:48.46" />
                    <SPLIT distance="1400" swimtime="00:18:28.03" />
                    <SPLIT distance="1450" swimtime="00:19:06.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="458" swimtime="00:02:44.70" resultid="8369" heatid="10763" lane="6" entrytime="00:02:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:18.62" />
                    <SPLIT distance="150" swimtime="00:02:02.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="528" swimtime="00:01:10.67" resultid="8370" heatid="10819" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="450" swimtime="00:02:13.09" resultid="8371" heatid="10865" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:04.56" />
                    <SPLIT distance="150" swimtime="00:01:39.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="462" swimtime="00:04:44.54" resultid="8372" heatid="10944" lane="4" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:07.16" />
                    <SPLIT distance="150" swimtime="00:01:42.84" />
                    <SPLIT distance="200" swimtime="00:02:18.91" />
                    <SPLIT distance="250" swimtime="00:02:55.09" />
                    <SPLIT distance="300" swimtime="00:03:31.96" />
                    <SPLIT distance="350" swimtime="00:04:09.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-06" firstname="Andrzej" gender="M" lastname="Szufarski" nation="POL" athleteid="3981">
              <RESULTS>
                <RESULT eventid="1190" points="105" swimtime="00:04:01.51" resultid="8380" heatid="10720" lane="6" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.84" />
                    <SPLIT distance="100" swimtime="00:01:51.37" />
                    <SPLIT distance="150" swimtime="00:02:58.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="91" swimtime="00:00:53.38" resultid="8381" heatid="10742" lane="1" entrytime="00:00:54.00" />
                <RESULT eventid="1422" points="113" swimtime="00:00:46.30" resultid="8382" heatid="10827" lane="1" entrytime="00:00:46.00" />
                <RESULT eventid="1452" points="79" swimtime="00:02:00.42" resultid="8383" heatid="10845" lane="9" entrytime="00:01:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="136" swimtime="00:00:51.27" resultid="8384" heatid="10914" lane="9" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="3959">
              <RESULTS>
                <RESULT eventid="1128" points="226" swimtime="00:23:48.65" resultid="8361" heatid="10677" lane="8" entrytime="00:23:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="100" swimtime="00:01:24.84" />
                    <SPLIT distance="150" swimtime="00:02:11.45" />
                    <SPLIT distance="200" swimtime="00:02:58.50" />
                    <SPLIT distance="250" swimtime="00:03:46.11" />
                    <SPLIT distance="300" swimtime="00:04:33.22" />
                    <SPLIT distance="350" swimtime="00:05:21.03" />
                    <SPLIT distance="400" swimtime="00:06:08.92" />
                    <SPLIT distance="450" swimtime="00:06:57.41" />
                    <SPLIT distance="500" swimtime="00:07:46.07" />
                    <SPLIT distance="550" swimtime="00:08:34.50" />
                    <SPLIT distance="600" swimtime="00:09:23.06" />
                    <SPLIT distance="650" swimtime="00:10:11.61" />
                    <SPLIT distance="700" swimtime="00:10:59.83" />
                    <SPLIT distance="750" swimtime="00:11:48.31" />
                    <SPLIT distance="800" swimtime="00:12:36.60" />
                    <SPLIT distance="850" swimtime="00:13:24.95" />
                    <SPLIT distance="900" swimtime="00:14:13.16" />
                    <SPLIT distance="950" swimtime="00:15:01.93" />
                    <SPLIT distance="1000" swimtime="00:15:50.44" />
                    <SPLIT distance="1050" swimtime="00:16:33.68" />
                    <SPLIT distance="1100" swimtime="00:17:27.12" />
                    <SPLIT distance="1150" swimtime="00:18:15.56" />
                    <SPLIT distance="1200" swimtime="00:19:03.17" />
                    <SPLIT distance="1250" swimtime="00:19:51.23" />
                    <SPLIT distance="1300" swimtime="00:20:39.06" />
                    <SPLIT distance="1350" swimtime="00:21:27.54" />
                    <SPLIT distance="1400" swimtime="00:22:15.12" />
                    <SPLIT distance="1450" swimtime="00:23:02.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="215" swimtime="00:03:10.01" resultid="8362" heatid="10723" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="100" swimtime="00:01:30.16" />
                    <SPLIT distance="150" swimtime="00:02:26.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="288" swimtime="00:01:11.00" resultid="8363" heatid="10778" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="301" swimtime="00:00:33.46" resultid="8364" heatid="10830" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1482" points="217" swimtime="00:02:49.66" resultid="8365" heatid="10860" lane="1" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:20.67" />
                    <SPLIT distance="150" swimtime="00:02:05.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="8366" heatid="10888" lane="9" entrytime="00:01:21.00" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="8367" heatid="10940" lane="3" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="3940">
              <RESULTS>
                <RESULT eventid="1160" points="122" swimtime="00:00:42.05" resultid="8345" heatid="10692" lane="0" entrytime="00:00:43.50" />
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="8346" heatid="10741" lane="0" entrytime="00:01:06.60" />
                <RESULT eventid="1452" points="50" swimtime="00:02:20.29" resultid="8347" heatid="10844" lane="0" entrytime="00:02:20.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="62" swimtime="00:04:17.40" resultid="8348" heatid="10857" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.18" />
                    <SPLIT distance="100" swimtime="00:01:54.49" />
                    <SPLIT distance="150" swimtime="00:03:04.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="39" swimtime="00:05:28.25" resultid="8349" heatid="10899" lane="3" entrytime="00:04:58.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.16" />
                    <SPLIT distance="100" swimtime="00:02:45.29" />
                    <SPLIT distance="150" swimtime="00:04:09.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-06" firstname="Arkadiusz" gender="M" lastname="Doliński" nation="POL" athleteid="3931">
              <RESULTS>
                <RESULT eventid="1098" points="186" swimtime="00:13:11.19" resultid="8337" heatid="10668" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:20.31" />
                    <SPLIT distance="150" swimtime="00:01:51.28" />
                    <SPLIT distance="200" swimtime="00:02:53.91" />
                    <SPLIT distance="250" swimtime="00:03:43.39" />
                    <SPLIT distance="300" swimtime="00:04:34.08" />
                    <SPLIT distance="350" swimtime="00:05:25.25" />
                    <SPLIT distance="400" swimtime="00:06:16.66" />
                    <SPLIT distance="450" swimtime="00:07:08.64" />
                    <SPLIT distance="500" swimtime="00:08:01.37" />
                    <SPLIT distance="550" swimtime="00:08:53.70" />
                    <SPLIT distance="600" swimtime="00:09:46.32" />
                    <SPLIT distance="650" swimtime="00:10:38.09" />
                    <SPLIT distance="700" swimtime="00:11:29.96" />
                    <SPLIT distance="750" swimtime="00:12:21.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="248" swimtime="00:03:01.38" resultid="8338" heatid="10719" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:21.72" />
                    <SPLIT distance="150" swimtime="00:02:18.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="327" swimtime="00:00:34.89" resultid="8339" heatid="10740" lane="1" />
                <RESULT eventid="1332" points="168" swimtime="00:03:21.80" resultid="8340" heatid="10791" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                    <SPLIT distance="100" swimtime="00:01:33.99" />
                    <SPLIT distance="150" swimtime="00:02:28.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="278" swimtime="00:01:19.42" resultid="8341" heatid="10843" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="228" swimtime="00:02:46.73" resultid="8342" heatid="10856" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:17.08" />
                    <SPLIT distance="150" swimtime="00:02:02.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="237" swimtime="00:03:00.61" resultid="8343" heatid="10899" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:25.59" />
                    <SPLIT distance="150" swimtime="00:02:14.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="8344" heatid="10935" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-25" firstname="Katarzyna" gender="F" lastname="Walenta" nation="POL" athleteid="3973">
              <RESULTS>
                <RESULT eventid="1144" points="515" swimtime="00:00:29.59" resultid="8373" heatid="10680" lane="5" />
                <RESULT eventid="1175" points="466" swimtime="00:02:42.64" resultid="8374" heatid="10718" lane="8" entrytime="00:02:44.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:02:04.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="421" swimtime="00:03:05.55" resultid="8375" heatid="10756" lane="2" entrytime="00:03:01.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:01:29.41" />
                    <SPLIT distance="150" swimtime="00:02:17.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="426" swimtime="00:01:25.49" resultid="8376" heatid="10808" lane="8" entrytime="00:01:25.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="416" swimtime="00:05:56.65" resultid="8377" heatid="10875" lane="6" entrytime="00:05:55.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="100" swimtime="00:01:24.04" />
                    <SPLIT distance="150" swimtime="00:02:10.76" />
                    <SPLIT distance="200" swimtime="00:02:56.49" />
                    <SPLIT distance="250" swimtime="00:03:45.39" />
                    <SPLIT distance="300" swimtime="00:04:34.43" />
                    <SPLIT distance="350" swimtime="00:05:16.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="407" swimtime="00:00:39.77" resultid="8378" heatid="10910" lane="3" entrytime="00:00:39.40" />
                <RESULT eventid="1674" points="386" swimtime="00:05:24.60" resultid="8379" heatid="10934" lane="0" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:17.64" />
                    <SPLIT distance="150" swimtime="00:01:59.17" />
                    <SPLIT distance="200" swimtime="00:02:41.15" />
                    <SPLIT distance="250" swimtime="00:03:22.77" />
                    <SPLIT distance="300" swimtime="00:04:04.14" />
                    <SPLIT distance="350" swimtime="00:04:44.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1518" points="73" swimtime="00:03:22.64" resultid="8385" heatid="10870" lane="0" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.66" />
                    <SPLIT distance="100" swimtime="00:01:30.88" />
                    <SPLIT distance="150" swimtime="00:02:09.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3951" number="1" />
                    <RELAYPOSITION athleteid="3946" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3940" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3981" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1368" points="48" swimtime="00:04:16.80" resultid="8386" heatid="10800" lane="0" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.66" />
                    <SPLIT distance="150" swimtime="00:01:30.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3951" number="1" />
                    <RELAYPOSITION athleteid="3946" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3981" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3940" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1518" status="DNS" swimtime="00:00:00.00" resultid="8387" heatid="10871" lane="6" entrytime="00:01:58.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3959" number="1" />
                    <RELAYPOSITION athleteid="3924" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3931" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3967" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1368" points="335" swimtime="00:02:14.47" resultid="8388" heatid="10801" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:08.77" />
                    <SPLIT distance="150" swimtime="00:01:42.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3931" number="1" />
                    <RELAYPOSITION athleteid="3967" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3959" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3924" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TRTOR" nation="POL" region="KUJ" clubid="3505" name="Toruński Klub Triathlonowy">
          <CONTACT city="Toruń" email="agusianamberone@poczta.onet.pl" name="Kostyra Agnieszka" phone="722053277" state="KUJ" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-16" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="3506">
              <RESULTS>
                <RESULT eventid="1113" points="228" swimtime="00:25:14.89" resultid="3507" heatid="10674" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                    <SPLIT distance="100" swimtime="00:01:35.97" />
                    <SPLIT distance="150" swimtime="00:02:27.43" />
                    <SPLIT distance="200" swimtime="00:03:19.51" />
                    <SPLIT distance="250" swimtime="00:04:11.40" />
                    <SPLIT distance="300" swimtime="00:05:03.39" />
                    <SPLIT distance="350" swimtime="00:05:54.02" />
                    <SPLIT distance="400" swimtime="00:06:45.96" />
                    <SPLIT distance="450" swimtime="00:07:37.06" />
                    <SPLIT distance="500" swimtime="00:08:28.08" />
                    <SPLIT distance="550" swimtime="00:09:17.78" />
                    <SPLIT distance="600" swimtime="00:10:08.52" />
                    <SPLIT distance="650" swimtime="00:10:58.79" />
                    <SPLIT distance="700" swimtime="00:11:50.31" />
                    <SPLIT distance="750" swimtime="00:12:40.37" />
                    <SPLIT distance="800" swimtime="00:13:31.19" />
                    <SPLIT distance="850" swimtime="00:14:21.35" />
                    <SPLIT distance="900" swimtime="00:15:12.29" />
                    <SPLIT distance="950" swimtime="00:16:02.47" />
                    <SPLIT distance="1000" swimtime="00:16:53.11" />
                    <SPLIT distance="1050" swimtime="00:17:43.13" />
                    <SPLIT distance="1100" swimtime="00:18:34.49" />
                    <SPLIT distance="1150" swimtime="00:19:24.49" />
                    <SPLIT distance="1200" swimtime="00:20:15.15" />
                    <SPLIT distance="1250" swimtime="00:21:06.00" />
                    <SPLIT distance="1300" swimtime="00:21:57.66" />
                    <SPLIT distance="1350" swimtime="00:22:47.83" />
                    <SPLIT distance="1400" swimtime="00:23:38.92" />
                    <SPLIT distance="1450" swimtime="00:24:27.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="394" swimtime="00:00:32.36" resultid="3508" heatid="10685" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1175" points="321" swimtime="00:03:04.17" resultid="3509" heatid="10716" lane="7" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                    <SPLIT distance="100" swimtime="00:01:28.25" />
                    <SPLIT distance="150" swimtime="00:02:20.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="266" swimtime="00:03:36.14" resultid="3510" heatid="10756" lane="8" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.11" />
                    <SPLIT distance="100" swimtime="00:01:43.94" />
                    <SPLIT distance="150" swimtime="00:02:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1317" points="149" swimtime="00:03:49.70" resultid="3511" heatid="10790" lane="0" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                    <SPLIT distance="100" swimtime="00:01:44.23" />
                    <SPLIT distance="150" swimtime="00:02:48.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="292" swimtime="00:02:50.27" resultid="3512" heatid="10854" lane="4" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:18.23" />
                    <SPLIT distance="150" swimtime="00:02:03.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="277" swimtime="00:06:48.51" resultid="3513" heatid="10875" lane="9" entrytime="00:06:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                    <SPLIT distance="100" swimtime="00:01:42.26" />
                    <SPLIT distance="150" swimtime="00:02:33.21" />
                    <SPLIT distance="200" swimtime="00:03:22.24" />
                    <SPLIT distance="250" swimtime="00:04:16.85" />
                    <SPLIT distance="300" swimtime="00:05:12.90" />
                    <SPLIT distance="350" swimtime="00:06:01.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="288" swimtime="00:03:07.65" resultid="3514" heatid="10896" lane="6" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.70" />
                    <SPLIT distance="100" swimtime="00:01:32.32" />
                    <SPLIT distance="150" swimtime="00:02:20.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="266" swimtime="00:06:07.36" resultid="3515" heatid="10933" lane="0" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:01:27.56" />
                    <SPLIT distance="150" swimtime="00:02:14.56" />
                    <SPLIT distance="200" swimtime="00:03:01.81" />
                    <SPLIT distance="250" swimtime="00:03:49.61" />
                    <SPLIT distance="300" swimtime="00:04:37.90" />
                    <SPLIT distance="350" swimtime="00:05:24.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-06-08" firstname="Mateusz" gender="M" lastname="Pałczyński" nation="POL" athleteid="3516">
              <RESULTS>
                <RESULT eventid="1098" points="221" swimtime="00:12:27.08" resultid="3517" heatid="10671" lane="7" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:01:59.93" />
                    <SPLIT distance="200" swimtime="00:02:44.05" />
                    <SPLIT distance="250" swimtime="00:03:28.85" />
                    <SPLIT distance="300" swimtime="00:04:15.46" />
                    <SPLIT distance="350" swimtime="00:05:03.61" />
                    <SPLIT distance="400" swimtime="00:05:52.03" />
                    <SPLIT distance="450" swimtime="00:06:41.11" />
                    <SPLIT distance="500" swimtime="00:07:30.71" />
                    <SPLIT distance="550" swimtime="00:08:19.34" />
                    <SPLIT distance="600" swimtime="00:09:09.51" />
                    <SPLIT distance="650" swimtime="00:09:59.55" />
                    <SPLIT distance="700" swimtime="00:10:49.51" />
                    <SPLIT distance="750" swimtime="00:11:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="383" swimtime="00:00:28.77" resultid="3518" heatid="10707" lane="8" entrytime="00:00:27.05" />
                <RESULT eventid="1190" points="371" swimtime="00:02:38.53" resultid="3519" heatid="10728" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                    <SPLIT distance="150" swimtime="00:01:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="338" swimtime="00:03:02.22" resultid="3520" heatid="10763" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:01:26.52" />
                    <SPLIT distance="150" swimtime="00:02:15.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="216" swimtime="00:03:05.59" resultid="3521" heatid="10794" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:22.33" />
                    <SPLIT distance="150" swimtime="00:02:12.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="416" swimtime="00:01:16.50" resultid="3522" heatid="10819" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="310" swimtime="00:06:00.11" resultid="3523" heatid="10880" lane="9" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:02:04.51" />
                    <SPLIT distance="200" swimtime="00:02:51.10" />
                    <SPLIT distance="250" swimtime="00:03:41.61" />
                    <SPLIT distance="300" swimtime="00:04:33.72" />
                    <SPLIT distance="350" swimtime="00:05:17.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="225" swimtime="00:03:03.95" resultid="3524" heatid="10902" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                    <SPLIT distance="100" swimtime="00:01:28.55" />
                    <SPLIT distance="150" swimtime="00:02:15.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="478" swimtime="00:00:33.77" resultid="3525" heatid="10925" lane="2" entrytime="00:00:32.45" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" nation="POL" region="WIE" clubid="4556" name="TS Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="4557">
              <RESULTS>
                <RESULT eventid="1098" points="190" swimtime="00:13:06.22" resultid="4558" heatid="10670" lane="6" entrytime="00:12:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                    <SPLIT distance="100" swimtime="00:01:31.95" />
                    <SPLIT distance="150" swimtime="00:02:21.50" />
                    <SPLIT distance="200" swimtime="00:03:12.19" />
                    <SPLIT distance="250" swimtime="00:04:02.34" />
                    <SPLIT distance="300" swimtime="00:04:52.47" />
                    <SPLIT distance="350" swimtime="00:05:42.69" />
                    <SPLIT distance="400" swimtime="00:06:33.05" />
                    <SPLIT distance="450" swimtime="00:07:22.94" />
                    <SPLIT distance="500" swimtime="00:08:12.62" />
                    <SPLIT distance="550" swimtime="00:09:01.37" />
                    <SPLIT distance="600" swimtime="00:09:50.98" />
                    <SPLIT distance="650" swimtime="00:10:39.73" />
                    <SPLIT distance="700" swimtime="00:11:29.31" />
                    <SPLIT distance="750" swimtime="00:12:18.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="203" swimtime="00:03:13.67" resultid="4559" heatid="10722" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                    <SPLIT distance="100" swimtime="00:01:35.96" />
                    <SPLIT distance="150" swimtime="00:02:30.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="164" swimtime="00:00:43.86" resultid="4560" heatid="10745" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="1332" status="DNS" swimtime="00:00:00.00" resultid="4561" heatid="10793" lane="9" entrytime="00:03:45.00" />
                <RESULT eventid="1452" points="182" swimtime="00:01:31.46" resultid="4562" heatid="10846" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="204" swimtime="00:06:53.93" resultid="4563" heatid="10878" lane="1" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.70" />
                    <SPLIT distance="100" swimtime="00:01:47.65" />
                    <SPLIT distance="150" swimtime="00:02:39.22" />
                    <SPLIT distance="200" swimtime="00:03:29.98" />
                    <SPLIT distance="250" swimtime="00:04:26.07" />
                    <SPLIT distance="300" swimtime="00:05:22.83" />
                    <SPLIT distance="350" swimtime="00:06:09.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="174" swimtime="00:03:20.17" resultid="4564" heatid="10901" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.38" />
                    <SPLIT distance="100" swimtime="00:01:37.92" />
                    <SPLIT distance="150" swimtime="00:02:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="183" swimtime="00:06:27.53" resultid="4565" heatid="10939" lane="7" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                    <SPLIT distance="100" swimtime="00:01:30.84" />
                    <SPLIT distance="150" swimtime="00:02:20.07" />
                    <SPLIT distance="200" swimtime="00:03:09.76" />
                    <SPLIT distance="250" swimtime="00:03:59.47" />
                    <SPLIT distance="300" swimtime="00:04:49.90" />
                    <SPLIT distance="350" swimtime="00:05:39.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="4575">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat I 65-69 lat" eventid="1059" points="163" swimtime="00:14:46.65" resultid="4576" heatid="10666" lane="3" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.80" />
                    <SPLIT distance="100" swimtime="00:01:46.76" />
                    <SPLIT distance="150" swimtime="00:02:43.98" />
                    <SPLIT distance="200" swimtime="00:03:41.24" />
                    <SPLIT distance="250" swimtime="00:04:38.32" />
                    <SPLIT distance="300" swimtime="00:05:35.10" />
                    <SPLIT distance="350" swimtime="00:06:31.75" />
                    <SPLIT distance="400" swimtime="00:07:26.28" />
                    <SPLIT distance="450" swimtime="00:08:22.16" />
                    <SPLIT distance="500" swimtime="00:09:18.20" />
                    <SPLIT distance="550" swimtime="00:10:14.76" />
                    <SPLIT distance="600" swimtime="00:11:10.90" />
                    <SPLIT distance="650" swimtime="00:12:05.63" />
                    <SPLIT distance="700" swimtime="00:13:00.78" />
                    <SPLIT distance="750" swimtime="00:13:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="215" swimtime="00:00:39.59" resultid="4577" heatid="10683" lane="9" entrytime="00:00:42.00" />
                <RESULT eventid="1226" points="158" swimtime="00:00:49.95" resultid="4578" heatid="10735" lane="3" entrytime="00:00:51.00" />
                <RESULT eventid="1287" points="166" swimtime="00:01:34.62" resultid="4579" heatid="10766" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="123" swimtime="00:00:49.06" resultid="4580" heatid="10821" lane="0" entrytime="00:00:51.00" />
                <RESULT eventid="1467" points="157" swimtime="00:03:29.03" resultid="4581" heatid="10852" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.65" />
                    <SPLIT distance="100" swimtime="00:01:44.94" />
                    <SPLIT distance="150" swimtime="00:02:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="163" swimtime="00:00:53.96" resultid="4582" heatid="10906" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="1674" points="152" swimtime="00:07:22.98" resultid="4583" heatid="10931" lane="3" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                    <SPLIT distance="100" swimtime="00:01:46.94" />
                    <SPLIT distance="150" swimtime="00:02:44.79" />
                    <SPLIT distance="200" swimtime="00:03:42.34" />
                    <SPLIT distance="250" swimtime="00:04:36.93" />
                    <SPLIT distance="300" swimtime="00:05:32.95" />
                    <SPLIT distance="350" swimtime="00:06:28.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Jacek" gender="M" lastname="Matyszczak" nation="POL" athleteid="4566">
              <RESULTS>
                <RESULT eventid="1160" points="419" swimtime="00:00:27.93" resultid="4567" heatid="10704" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="1190" points="273" swimtime="00:02:55.53" resultid="4568" heatid="10724" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:02:15.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="241" swimtime="00:00:38.63" resultid="4569" heatid="10746" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="1302" points="395" swimtime="00:01:03.89" resultid="4570" heatid="10783" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="347" swimtime="00:00:31.90" resultid="4571" heatid="10831" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1482" points="298" swimtime="00:02:32.62" resultid="4572" heatid="10861" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:12.53" />
                    <SPLIT distance="150" swimtime="00:01:53.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="183" swimtime="00:03:16.80" resultid="4573" heatid="10901" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.35" />
                    <SPLIT distance="100" swimtime="00:01:35.79" />
                    <SPLIT distance="150" swimtime="00:02:27.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="278" swimtime="00:05:36.89" resultid="4574" heatid="10941" lane="5" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                    <SPLIT distance="100" swimtime="00:01:14.01" />
                    <SPLIT distance="150" swimtime="00:01:55.68" />
                    <SPLIT distance="200" swimtime="00:02:38.94" />
                    <SPLIT distance="250" swimtime="00:03:23.08" />
                    <SPLIT distance="300" swimtime="00:04:08.19" />
                    <SPLIT distance="350" swimtime="00:04:53.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BULOM" nation="POL" region="PDL" clubid="3367" name="UKS Butterfly">
          <CONTACT city="Łomża" email="jarekszeremet@wp.pl" name="Szeremet Jarosław" phone="502277492" state="PDL" street="Rycerska /73" zip="18-400" />
          <ATHLETES>
            <ATHLETE birthdate="1986-03-16" firstname="Bartosz" gender="M" lastname="Kutny" nation="POL" license="101009700023" athleteid="3368">
              <RESULTS>
                <RESULT eventid="1128" points="304" swimtime="00:21:34.80" resultid="6954" heatid="10678" lane="5" entrytime="00:21:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:09.80" />
                    <SPLIT distance="150" swimtime="00:01:49.66" />
                    <SPLIT distance="200" swimtime="00:02:30.35" />
                    <SPLIT distance="250" swimtime="00:03:12.22" />
                    <SPLIT distance="300" swimtime="00:03:54.61" />
                    <SPLIT distance="350" swimtime="00:04:37.22" />
                    <SPLIT distance="400" swimtime="00:05:20.17" />
                    <SPLIT distance="450" swimtime="00:06:04.10" />
                    <SPLIT distance="500" swimtime="00:06:48.13" />
                    <SPLIT distance="550" swimtime="00:07:32.44" />
                    <SPLIT distance="600" swimtime="00:08:16.54" />
                    <SPLIT distance="650" swimtime="00:09:01.35" />
                    <SPLIT distance="700" swimtime="00:09:45.56" />
                    <SPLIT distance="750" swimtime="00:10:30.43" />
                    <SPLIT distance="800" swimtime="00:11:14.47" />
                    <SPLIT distance="850" swimtime="00:11:59.21" />
                    <SPLIT distance="900" swimtime="00:12:43.61" />
                    <SPLIT distance="950" swimtime="00:13:28.63" />
                    <SPLIT distance="1000" swimtime="00:14:13.24" />
                    <SPLIT distance="1050" swimtime="00:14:57.85" />
                    <SPLIT distance="1100" swimtime="00:15:42.68" />
                    <SPLIT distance="1150" swimtime="00:16:27.58" />
                    <SPLIT distance="1200" swimtime="00:17:12.63" />
                    <SPLIT distance="1250" swimtime="00:17:57.80" />
                    <SPLIT distance="1300" swimtime="00:18:42.75" />
                    <SPLIT distance="1350" swimtime="00:19:26.84" />
                    <SPLIT distance="1400" swimtime="00:20:10.64" />
                    <SPLIT distance="1450" swimtime="00:20:54.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="418" swimtime="00:00:27.95" resultid="6955" heatid="10706" lane="7" entrytime="00:00:27.50" entrycourse="SCM" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="6956" heatid="10725" lane="5" entrytime="00:02:48.00" entrycourse="SCM" />
                <RESULT eventid="1242" points="326" swimtime="00:00:34.90" resultid="6957" heatid="10745" lane="8" entrytime="00:00:40.01" entrycourse="SCM" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="6958" heatid="10783" lane="0" entrytime="00:01:03.00" entrycourse="SCM" />
                <RESULT eventid="1422" points="380" swimtime="00:00:30.95" resultid="6959" heatid="10834" lane="2" entrytime="00:00:30.01" entrycourse="SCM" />
                <RESULT eventid="1482" points="350" swimtime="00:02:24.73" resultid="6960" heatid="10862" lane="2" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                    <SPLIT distance="150" swimtime="00:01:47.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" status="DNS" swimtime="00:00:00.00" resultid="6961" heatid="10881" lane="2" entrytime="00:05:10.00" entrycourse="SCM" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="6962" heatid="10888" lane="7" entrytime="00:01:18.00" entrycourse="SCM" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="6963" heatid="10918" lane="8" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CIPOZ" nation="POL" region="WLK" clubid="4584" name="UKS CITYZEN Poznań">
          <CONTACT city="Poznań" email="oskar.borowczyk@gmail.com" name="Borowczyk" phone="730979848" street="Droga Dębińska" zip="60-555" />
          <ATHLETES>
            <ATHLETE birthdate="1974-08-05" firstname="Kinga" gender="F" lastname="Jaruga" nation="POL" athleteid="4585">
              <RESULTS>
                <RESULT eventid="1059" points="259" swimtime="00:12:40.34" resultid="7901" heatid="10667" lane="6" entrytime="00:12:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                    <SPLIT distance="100" swimtime="00:01:26.19" />
                    <SPLIT distance="150" swimtime="00:02:13.03" />
                    <SPLIT distance="200" swimtime="00:03:00.70" />
                    <SPLIT distance="250" swimtime="00:03:48.59" />
                    <SPLIT distance="300" swimtime="00:04:36.47" />
                    <SPLIT distance="350" swimtime="00:05:24.75" />
                    <SPLIT distance="400" swimtime="00:06:13.18" />
                    <SPLIT distance="450" swimtime="00:07:01.89" />
                    <SPLIT distance="500" swimtime="00:07:51.20" />
                    <SPLIT distance="550" swimtime="00:08:40.44" />
                    <SPLIT distance="600" swimtime="00:09:29.27" />
                    <SPLIT distance="650" swimtime="00:10:17.94" />
                    <SPLIT distance="700" swimtime="00:11:06.04" />
                    <SPLIT distance="750" swimtime="00:11:54.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="298" swimtime="00:01:17.94" resultid="7902" heatid="10768" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="257" swimtime="00:00:38.41" resultid="7903" heatid="10822" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="1467" points="286" swimtime="00:02:51.34" resultid="7904" heatid="10853" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:02:06.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="182" swimtime="00:01:37.77" resultid="7905" heatid="10883" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="270" swimtime="00:06:05.77" resultid="7906" heatid="10933" lane="6" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:24.13" />
                    <SPLIT distance="150" swimtime="00:02:10.74" />
                    <SPLIT distance="200" swimtime="00:02:58.07" />
                    <SPLIT distance="250" swimtime="00:03:45.80" />
                    <SPLIT distance="300" swimtime="00:04:33.50" />
                    <SPLIT distance="350" swimtime="00:05:20.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08314" nation="POL" region="14" clubid="4112" name="UKS Delfin Garwolin">
          <CONTACT city="Garwolin" email="uksdelfingarwolin@o2.pl" internet="www.uksdelfingarwolin.pl" name="Mianowski" phone="792843291" state="MAZOW" street="Olimpijska" zip="08-400" />
          <ATHLETES>
            <ATHLETE birthdate="1996-12-29" firstname="Mateusz" gender="M" lastname="Szczypek" nation="POL" athleteid="4113">
              <RESULTS>
                <RESULT eventid="1098" points="314" swimtime="00:11:04.57" resultid="6472" heatid="10671" lane="4" entrytime="00:11:24.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:11.65" />
                    <SPLIT distance="150" swimtime="00:01:51.50" />
                    <SPLIT distance="200" swimtime="00:02:31.82" />
                    <SPLIT distance="250" swimtime="00:03:12.57" />
                    <SPLIT distance="300" swimtime="00:03:54.17" />
                    <SPLIT distance="350" swimtime="00:04:35.94" />
                    <SPLIT distance="400" swimtime="00:05:18.54" />
                    <SPLIT distance="450" swimtime="00:06:01.51" />
                    <SPLIT distance="500" swimtime="00:06:45.83" />
                    <SPLIT distance="550" swimtime="00:07:29.63" />
                    <SPLIT distance="600" swimtime="00:08:13.54" />
                    <SPLIT distance="650" swimtime="00:08:57.14" />
                    <SPLIT distance="700" swimtime="00:09:41.14" />
                    <SPLIT distance="750" swimtime="00:10:24.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="428" swimtime="00:00:27.74" resultid="6473" heatid="10706" lane="5" entrytime="00:00:27.47" />
                <RESULT eventid="1190" points="361" swimtime="00:02:40.00" resultid="6474" heatid="10727" lane="2" entrytime="00:02:38.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:02:01.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="435" swimtime="00:01:01.89" resultid="6475" heatid="10785" lane="9" entrytime="00:01:00.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="434" swimtime="00:00:29.61" resultid="6476" heatid="10835" lane="7" entrytime="00:00:29.60" />
                <RESULT eventid="1482" points="387" swimtime="00:02:19.95" resultid="6477" heatid="10863" lane="3" entrytime="00:02:18.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:07.02" />
                    <SPLIT distance="150" swimtime="00:01:44.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="482" swimtime="00:00:33.68" resultid="6478" heatid="10924" lane="3" entrytime="00:00:33.68" />
                <RESULT eventid="1695" points="353" swimtime="00:05:11.32" resultid="6479" heatid="10942" lane="7" entrytime="00:05:13.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:12.71" />
                    <SPLIT distance="150" swimtime="00:01:52.90" />
                    <SPLIT distance="200" swimtime="00:02:33.09" />
                    <SPLIT distance="250" swimtime="00:03:13.46" />
                    <SPLIT distance="300" swimtime="00:03:53.62" />
                    <SPLIT distance="350" swimtime="00:04:34.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" region="14" clubid="3341" name="Uks Delfin Legionowo">
          <CONTACT city="LEGIONOWO" email="delfin-trener@wp.pl" internet="www.delfinlegionowo.pl" name="RAFAŁ PERL" phone="601 436 700" state="MAZ" street="KRÓLOWEJ JADWIGI 11" zip="05-120" />
          <ATHLETES>
            <ATHLETE birthdate="1996-06-07" firstname="Michał" gender="M" lastname="Perl" nation="POL" athleteid="6844">
              <RESULTS>
                <RESULT eventid="1160" points="601" swimtime="00:00:24.77" resultid="6845" heatid="10711" lane="4" entrytime="00:00:23.57" />
                <RESULT eventid="1422" points="557" swimtime="00:00:27.25" resultid="6846" heatid="10837" lane="0" entrytime="00:00:28.02" />
                <RESULT eventid="1638" points="653" swimtime="00:00:30.44" resultid="6847" heatid="10926" lane="4" entrytime="00:00:28.95" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="PDK" clubid="4670" name="Uks Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1972-01-17" firstname="Sławomir" gender="M" lastname="Kowalski" nation="POL" athleteid="4682">
              <RESULTS>
                <RESULT eventid="1098" points="253" swimtime="00:11:54.70" resultid="8225" heatid="10670" lane="8" entrytime="00:13:22.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:17.59" />
                    <SPLIT distance="150" swimtime="00:02:01.00" />
                    <SPLIT distance="200" swimtime="00:02:45.68" />
                    <SPLIT distance="250" swimtime="00:03:30.31" />
                    <SPLIT distance="300" swimtime="00:04:16.04" />
                    <SPLIT distance="350" swimtime="00:05:02.11" />
                    <SPLIT distance="400" swimtime="00:05:48.76" />
                    <SPLIT distance="450" swimtime="00:06:34.95" />
                    <SPLIT distance="500" swimtime="00:07:22.13" />
                    <SPLIT distance="550" swimtime="00:08:08.53" />
                    <SPLIT distance="600" swimtime="00:08:55.77" />
                    <SPLIT distance="650" swimtime="00:09:41.76" />
                    <SPLIT distance="700" swimtime="00:10:28.57" />
                    <SPLIT distance="750" swimtime="00:11:13.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="376" swimtime="00:00:28.95" resultid="8226" heatid="10690" lane="2" />
                <RESULT eventid="1190" points="324" swimtime="00:02:45.96" resultid="8227" heatid="10725" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:19.09" />
                    <SPLIT distance="150" swimtime="00:02:06.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="343" swimtime="00:03:01.31" resultid="8228" heatid="10762" lane="8" entrytime="00:02:59.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                    <SPLIT distance="100" swimtime="00:01:28.39" />
                    <SPLIT distance="150" swimtime="00:02:15.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="380" swimtime="00:01:18.85" resultid="8229" heatid="10816" lane="7" entrytime="00:01:21.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="8230" heatid="10831" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1638" points="444" swimtime="00:00:34.62" resultid="8231" heatid="10921" lane="7" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-30" firstname="Angelika" gender="F" lastname="Rozmus" nation="POL" athleteid="4727">
              <RESULTS>
                <RESULT eventid="1144" points="361" swimtime="00:00:33.30" resultid="8264" heatid="10686" lane="6" entrytime="00:00:32.50" />
                <RESULT eventid="1175" points="319" swimtime="00:03:04.55" resultid="8265" heatid="10717" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:27.81" />
                    <SPLIT distance="150" swimtime="00:02:20.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="286" swimtime="00:00:41.05" resultid="8266" heatid="10738" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1257" points="296" swimtime="00:03:28.65" resultid="8267" heatid="10755" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                    <SPLIT distance="100" swimtime="00:01:41.05" />
                    <SPLIT distance="150" swimtime="00:02:36.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="295" swimtime="00:01:36.56" resultid="8268" heatid="10808" lane="9" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="282" swimtime="00:06:45.72" resultid="8269" heatid="10874" lane="2" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                    <SPLIT distance="100" swimtime="00:01:34.85" />
                    <SPLIT distance="150" swimtime="00:02:30.19" />
                    <SPLIT distance="200" swimtime="00:03:23.13" />
                    <SPLIT distance="250" swimtime="00:04:20.51" />
                    <SPLIT distance="300" swimtime="00:05:16.61" />
                    <SPLIT distance="350" swimtime="00:06:02.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="231" swimtime="00:01:30.37" resultid="8270" heatid="10883" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="295" swimtime="00:00:44.28" resultid="8271" heatid="10910" lane="9" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-15" firstname="Witold" gender="M" lastname="Flak" nation="POL" athleteid="4712">
              <RESULTS>
                <RESULT eventid="1160" points="381" swimtime="00:00:28.82" resultid="8251" heatid="10703" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1242" points="283" swimtime="00:00:36.59" resultid="8252" heatid="10746" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1272" points="259" swimtime="00:03:19.03" resultid="8253" heatid="10760" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:33.65" />
                    <SPLIT distance="150" swimtime="00:02:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="315" swimtime="00:01:23.93" resultid="8254" heatid="10815" lane="4" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="8255" heatid="10829" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1638" points="376" swimtime="00:00:36.60" resultid="8256" heatid="10919" lane="3" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-14" firstname="Maciej" gender="M" lastname="Kunicki" nation="POL" athleteid="4671">
              <RESULTS>
                <RESULT eventid="1160" points="320" swimtime="00:00:30.54" resultid="8216" heatid="10702" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1332" points="222" swimtime="00:03:03.94" resultid="8217" heatid="10794" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                    <SPLIT distance="100" swimtime="00:01:27.16" />
                    <SPLIT distance="150" swimtime="00:02:15.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="335" swimtime="00:00:32.27" resultid="8218" heatid="10832" lane="1" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-25" firstname="Artur" gender="M" lastname="Szklarz" nation="POL" athleteid="4706">
              <RESULTS>
                <RESULT eventid="1098" points="305" swimtime="00:11:11.37" resultid="8246" heatid="10672" lane="0" entrytime="00:11:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:15.18" />
                    <SPLIT distance="150" swimtime="00:01:55.85" />
                    <SPLIT distance="200" swimtime="00:02:37.14" />
                    <SPLIT distance="250" swimtime="00:03:18.18" />
                    <SPLIT distance="300" swimtime="00:03:59.83" />
                    <SPLIT distance="350" swimtime="00:04:41.25" />
                    <SPLIT distance="400" swimtime="00:05:23.39" />
                    <SPLIT distance="450" swimtime="00:06:05.10" />
                    <SPLIT distance="500" swimtime="00:06:47.75" />
                    <SPLIT distance="550" swimtime="00:07:30.35" />
                    <SPLIT distance="600" swimtime="00:08:13.90" />
                    <SPLIT distance="650" swimtime="00:08:57.54" />
                    <SPLIT distance="700" swimtime="00:09:42.61" />
                    <SPLIT distance="750" swimtime="00:10:27.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="374" swimtime="00:00:29.02" resultid="8247" heatid="10702" lane="2" entrytime="00:00:29.09" />
                <RESULT eventid="1302" points="414" swimtime="00:01:02.90" resultid="8248" heatid="10782" lane="6" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="356" swimtime="00:00:31.62" resultid="8249" heatid="10831" lane="4" entrytime="00:00:32.50" />
                <RESULT eventid="1638" points="401" swimtime="00:00:35.82" resultid="8250" heatid="10921" lane="5" entrytime="00:00:36.79" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="4719">
              <RESULTS>
                <RESULT eventid="1160" points="446" swimtime="00:00:27.36" resultid="8257" heatid="10702" lane="8" entrytime="00:00:29.34" />
                <RESULT eventid="1190" points="385" swimtime="00:02:36.68" resultid="8258" heatid="10726" lane="4" entrytime="00:02:40.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:13.90" />
                    <SPLIT distance="150" swimtime="00:02:01.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="461" swimtime="00:01:00.72" resultid="8259" heatid="10784" lane="8" entrytime="00:01:01.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="397" swimtime="00:01:17.68" resultid="8260" heatid="10816" lane="2" entrytime="00:01:21.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="420" swimtime="00:02:16.16" resultid="8261" heatid="10864" lane="5" entrytime="00:02:14.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:01:05.68" />
                    <SPLIT distance="150" swimtime="00:01:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="8262" heatid="10889" lane="6" entrytime="00:01:11.02" />
                <RESULT eventid="1638" points="444" swimtime="00:00:34.62" resultid="8263" heatid="10922" lane="9" entrytime="00:00:36.28" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-14" firstname="Piotr" gender="M" lastname="Darowski" nation="POL" athleteid="4690">
              <RESULTS>
                <RESULT eventid="1190" points="383" swimtime="00:02:36.86" resultid="8232" heatid="10728" lane="5" entrytime="00:02:33.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:13.43" />
                    <SPLIT distance="150" swimtime="00:01:57.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="408" swimtime="00:02:51.21" resultid="8233" heatid="10763" lane="4" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:18.81" />
                    <SPLIT distance="150" swimtime="00:02:04.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="384" swimtime="00:01:18.57" resultid="8234" heatid="10817" lane="0" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="355" swimtime="00:05:44.09" resultid="8235" heatid="10880" lane="7" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:15.29" />
                    <SPLIT distance="150" swimtime="00:02:02.96" />
                    <SPLIT distance="200" swimtime="00:02:50.37" />
                    <SPLIT distance="250" swimtime="00:03:35.98" />
                    <SPLIT distance="300" swimtime="00:04:22.91" />
                    <SPLIT distance="350" swimtime="00:05:03.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="305" swimtime="00:01:13.97" resultid="8236" heatid="10889" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="426" swimtime="00:00:35.09" resultid="8237" heatid="10923" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="4697">
              <RESULTS>
                <RESULT eventid="1128" points="253" swimtime="00:22:56.99" resultid="8238" heatid="10678" lane="0" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="150" swimtime="00:02:00.29" />
                    <SPLIT distance="200" swimtime="00:02:42.96" />
                    <SPLIT distance="250" swimtime="00:03:26.96" />
                    <SPLIT distance="300" swimtime="00:04:11.00" />
                    <SPLIT distance="350" swimtime="00:04:55.89" />
                    <SPLIT distance="400" swimtime="00:05:41.20" />
                    <SPLIT distance="450" swimtime="00:06:27.08" />
                    <SPLIT distance="500" swimtime="00:07:13.15" />
                    <SPLIT distance="550" swimtime="00:07:58.91" />
                    <SPLIT distance="600" swimtime="00:08:45.61" />
                    <SPLIT distance="650" swimtime="00:09:31.71" />
                    <SPLIT distance="700" swimtime="00:10:18.74" />
                    <SPLIT distance="750" swimtime="00:11:05.15" />
                    <SPLIT distance="800" swimtime="00:11:52.04" />
                    <SPLIT distance="850" swimtime="00:12:38.75" />
                    <SPLIT distance="900" swimtime="00:13:25.65" />
                    <SPLIT distance="950" swimtime="00:14:12.68" />
                    <SPLIT distance="1000" swimtime="00:15:00.46" />
                    <SPLIT distance="1050" swimtime="00:15:48.24" />
                    <SPLIT distance="1100" swimtime="00:16:36.59" />
                    <SPLIT distance="1150" swimtime="00:17:24.89" />
                    <SPLIT distance="1200" swimtime="00:18:13.21" />
                    <SPLIT distance="1250" swimtime="00:19:02.11" />
                    <SPLIT distance="1300" swimtime="00:19:50.59" />
                    <SPLIT distance="1350" swimtime="00:20:38.53" />
                    <SPLIT distance="1400" swimtime="00:21:26.38" />
                    <SPLIT distance="1450" swimtime="00:22:12.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="297" swimtime="00:00:31.33" resultid="8239" heatid="10701" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="1302" points="323" swimtime="00:01:08.31" resultid="8240" heatid="10780" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="183" swimtime="00:03:16.30" resultid="8241" heatid="10794" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                    <SPLIT distance="100" swimtime="00:01:35.60" />
                    <SPLIT distance="150" swimtime="00:02:27.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="280" swimtime="00:02:35.81" resultid="8242" heatid="10862" lane="0" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                    <SPLIT distance="150" swimtime="00:01:53.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="244" swimtime="00:06:29.88" resultid="8243" heatid="10878" lane="6" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:26.87" />
                    <SPLIT distance="150" swimtime="00:02:21.55" />
                    <SPLIT distance="200" swimtime="00:03:13.29" />
                    <SPLIT distance="250" swimtime="00:04:09.70" />
                    <SPLIT distance="300" swimtime="00:05:05.36" />
                    <SPLIT distance="350" swimtime="00:05:49.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="214" swimtime="00:03:06.84" resultid="8244" heatid="10899" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="150" swimtime="00:02:22.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="291" swimtime="00:05:31.75" resultid="8245" heatid="10942" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                    <SPLIT distance="150" swimtime="00:01:59.68" />
                    <SPLIT distance="200" swimtime="00:02:41.84" />
                    <SPLIT distance="250" swimtime="00:03:25.41" />
                    <SPLIT distance="300" swimtime="00:04:08.48" />
                    <SPLIT distance="350" swimtime="00:04:52.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-27" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" athleteid="4675">
              <RESULTS>
                <RESULT eventid="1128" points="307" swimtime="00:21:30.11" resultid="8219" heatid="10679" lane="6" entrytime="00:19:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:16.10" />
                    <SPLIT distance="150" swimtime="00:01:57.98" />
                    <SPLIT distance="200" swimtime="00:02:40.97" />
                    <SPLIT distance="250" swimtime="00:03:24.40" />
                    <SPLIT distance="300" swimtime="00:04:08.30" />
                    <SPLIT distance="350" swimtime="00:04:52.33" />
                    <SPLIT distance="400" swimtime="00:05:36.37" />
                    <SPLIT distance="450" swimtime="00:06:20.14" />
                    <SPLIT distance="500" swimtime="00:07:03.53" />
                    <SPLIT distance="550" swimtime="00:07:47.38" />
                    <SPLIT distance="600" swimtime="00:08:30.94" />
                    <SPLIT distance="650" swimtime="00:09:14.04" />
                    <SPLIT distance="700" swimtime="00:09:57.65" />
                    <SPLIT distance="750" swimtime="00:10:41.39" />
                    <SPLIT distance="800" swimtime="00:11:25.34" />
                    <SPLIT distance="850" swimtime="00:12:09.27" />
                    <SPLIT distance="900" swimtime="00:12:52.89" />
                    <SPLIT distance="950" swimtime="00:13:36.55" />
                    <SPLIT distance="1000" swimtime="00:14:20.30" />
                    <SPLIT distance="1050" swimtime="00:15:03.73" />
                    <SPLIT distance="1100" swimtime="00:15:47.25" />
                    <SPLIT distance="1150" swimtime="00:16:31.04" />
                    <SPLIT distance="1200" swimtime="00:17:14.52" />
                    <SPLIT distance="1250" swimtime="00:17:57.28" />
                    <SPLIT distance="1300" swimtime="00:18:40.48" />
                    <SPLIT distance="1350" swimtime="00:19:23.41" />
                    <SPLIT distance="1400" swimtime="00:20:06.44" />
                    <SPLIT distance="1450" swimtime="00:20:48.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="8220" heatid="10690" lane="8" />
                <RESULT eventid="1272" points="472" swimtime="00:02:43.09" resultid="8221" heatid="10764" lane="3" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:17.24" />
                    <SPLIT distance="150" swimtime="00:01:59.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="8222" heatid="10809" lane="8" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="8223" heatid="10926" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="8224" heatid="10943" lane="3" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="375" swimtime="00:02:09.50" resultid="8272" heatid="10801" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:42.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4706" number="1" />
                    <RELAYPOSITION athleteid="4690" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4682" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4719" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" points="420" swimtime="00:01:53.30" resultid="8274" heatid="10872" lane="0" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                    <SPLIT distance="100" swimtime="00:00:57.14" />
                    <SPLIT distance="150" swimtime="00:01:26.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4712" number="1" />
                    <RELAYPOSITION athleteid="4706" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4682" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4719" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="DOL" clubid="3585" name="UKS Energetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" internet="www.plywanie-zgorzelec.pl" name="Kondracki Łukasz" phone="693852488" state="DOL" street="Maratońska 2" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="3597">
              <RESULTS>
                <RESULT eventid="1098" points="85" swimtime="00:17:05.86" resultid="9029" heatid="10669" lane="3" entrytime="00:16:30.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.08" />
                    <SPLIT distance="100" swimtime="00:01:58.18" />
                    <SPLIT distance="150" swimtime="00:03:02.88" />
                    <SPLIT distance="200" swimtime="00:04:09.35" />
                    <SPLIT distance="250" swimtime="00:05:14.79" />
                    <SPLIT distance="300" swimtime="00:06:22.10" />
                    <SPLIT distance="350" swimtime="00:07:25.65" />
                    <SPLIT distance="400" swimtime="00:08:30.44" />
                    <SPLIT distance="450" swimtime="00:09:33.50" />
                    <SPLIT distance="500" swimtime="00:10:38.50" />
                    <SPLIT distance="550" swimtime="00:11:43.65" />
                    <SPLIT distance="600" swimtime="00:12:49.53" />
                    <SPLIT distance="650" swimtime="00:13:55.02" />
                    <SPLIT distance="700" swimtime="00:15:00.35" />
                    <SPLIT distance="750" swimtime="00:16:04.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="117" swimtime="00:00:42.71" resultid="9030" heatid="10691" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1190" points="81" swimtime="00:04:23.13" resultid="9031" heatid="10720" lane="2" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.97" />
                    <SPLIT distance="100" swimtime="00:02:08.43" />
                    <SPLIT distance="150" swimtime="00:03:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="100" swimtime="00:00:51.71" resultid="9032" heatid="10741" lane="4" entrytime="00:00:55.00" />
                <RESULT eventid="1332" points="50" swimtime="00:05:01.59" resultid="9033" heatid="10792" lane="1" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.12" />
                    <SPLIT distance="100" swimtime="00:02:25.73" />
                    <SPLIT distance="150" swimtime="00:03:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="95" swimtime="00:01:53.49" resultid="9034" heatid="10845" lane="0" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="84" swimtime="00:09:15.96" resultid="9035" heatid="10877" lane="9" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.05" />
                    <SPLIT distance="100" swimtime="00:02:23.15" />
                    <SPLIT distance="150" swimtime="00:03:30.08" />
                    <SPLIT distance="200" swimtime="00:04:33.76" />
                    <SPLIT distance="250" swimtime="00:05:55.48" />
                    <SPLIT distance="300" swimtime="00:07:16.85" />
                    <SPLIT distance="350" swimtime="00:08:18.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="92" swimtime="00:04:07.21" resultid="9036" heatid="10900" lane="8" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.78" />
                    <SPLIT distance="100" swimtime="00:02:03.85" />
                    <SPLIT distance="150" swimtime="00:03:06.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="88" swimtime="00:08:14.55" resultid="9037" heatid="10936" lane="5" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.07" />
                    <SPLIT distance="100" swimtime="00:01:52.46" />
                    <SPLIT distance="150" swimtime="00:02:54.26" />
                    <SPLIT distance="200" swimtime="00:03:58.80" />
                    <SPLIT distance="250" swimtime="00:05:02.95" />
                    <SPLIT distance="300" swimtime="00:06:08.24" />
                    <SPLIT distance="350" swimtime="00:07:14.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="09914" nation="POL" region="14" clubid="9222" name="UKS Fala Nieporęt">
          <CONTACT name="Krawczak" phone="530077078" />
          <ATHLETES>
            <ATHLETE birthdate="1986-05-14" firstname="Bartosz" gender="M" lastname="Krawczak" nation="POL" athleteid="9223">
              <RESULTS>
                <RESULT eventid="1160" points="599" swimtime="00:00:24.80" resultid="9224" heatid="10711" lane="7" entrytime="00:00:24.50" />
                <RESULT eventid="1302" points="624" swimtime="00:00:54.87" resultid="9225" heatid="10788" lane="0" entrytime="00:00:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="9226" heatid="10837" lane="5" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="026" nation="POL" region="PDK" clubid="6061" name="UKS FREGATA Kolbuszowa">
          <CONTACT name="Pietryka" phone="604620876" />
          <ATHLETES>
            <ATHLETE birthdate="1986-07-20" firstname="Bartosz" gender="M" lastname="Pietryka" nation="POL" license="102608700019" athleteid="6062">
              <RESULTS>
                <RESULT eventid="1242" points="479" swimtime="00:00:30.71" resultid="6558" heatid="10750" lane="4" entrytime="00:00:30.20" entrycourse="LCM" />
                <RESULT eventid="1422" points="551" swimtime="00:00:27.35" resultid="6559" heatid="10837" lane="6" entrytime="00:00:27.50" entrycourse="LCM" />
                <RESULT eventid="1452" points="399" swimtime="00:01:10.38" resultid="6560" heatid="10850" lane="0" entrytime="00:01:06.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="550" swimtime="00:01:00.79" resultid="6561" heatid="10892" lane="0" entrytime="00:01:00.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="6562" heatid="10944" lane="7" entrytime="00:04:50.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="07614" nation="POL" region="14" clubid="5212" name="UKS GOS Raszyn">
          <CONTACT name="s" />
          <ATHLETES>
            <ATHLETE birthdate="1962-12-05" firstname="Leszek" gender="M" lastname="Rąpałą" nation="POL" athleteid="5213">
              <RESULTS>
                <RESULT eventid="1128" points="138" swimtime="00:28:02.17" resultid="7940" heatid="10675" lane="1" entrytime="00:29:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                    <SPLIT distance="100" swimtime="00:01:42.22" />
                    <SPLIT distance="150" swimtime="00:02:36.52" />
                    <SPLIT distance="200" swimtime="00:03:30.84" />
                    <SPLIT distance="250" swimtime="00:04:27.88" />
                    <SPLIT distance="300" swimtime="00:05:24.65" />
                    <SPLIT distance="350" swimtime="00:06:20.51" />
                    <SPLIT distance="400" swimtime="00:07:16.98" />
                    <SPLIT distance="450" swimtime="00:08:14.43" />
                    <SPLIT distance="500" swimtime="00:09:10.62" />
                    <SPLIT distance="550" swimtime="00:10:07.28" />
                    <SPLIT distance="600" swimtime="00:11:04.81" />
                    <SPLIT distance="650" swimtime="00:12:02.71" />
                    <SPLIT distance="700" swimtime="00:13:00.28" />
                    <SPLIT distance="750" swimtime="00:13:56.28" />
                    <SPLIT distance="800" swimtime="00:14:53.37" />
                    <SPLIT distance="850" swimtime="00:15:50.18" />
                    <SPLIT distance="900" swimtime="00:16:47.80" />
                    <SPLIT distance="950" swimtime="00:17:45.65" />
                    <SPLIT distance="1000" swimtime="00:18:43.75" />
                    <SPLIT distance="1050" swimtime="00:19:39.94" />
                    <SPLIT distance="1100" swimtime="00:20:36.70" />
                    <SPLIT distance="1150" swimtime="00:21:33.20" />
                    <SPLIT distance="1200" swimtime="00:22:29.46" />
                    <SPLIT distance="1250" swimtime="00:23:25.10" />
                    <SPLIT distance="1300" swimtime="00:24:22.86" />
                    <SPLIT distance="1350" swimtime="00:25:18.29" />
                    <SPLIT distance="1400" swimtime="00:26:13.32" />
                    <SPLIT distance="1450" swimtime="00:27:08.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="110" swimtime="00:03:57.51" resultid="7941" heatid="10720" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.92" />
                    <SPLIT distance="100" swimtime="00:02:00.77" />
                    <SPLIT distance="150" swimtime="00:03:08.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="106" swimtime="00:00:47.27" resultid="7942" heatid="10827" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1695" points="162" swimtime="00:06:43.55" resultid="7943" heatid="10937" lane="8" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.50" />
                    <SPLIT distance="100" swimtime="00:01:33.57" />
                    <SPLIT distance="150" swimtime="00:02:26.01" />
                    <SPLIT distance="200" swimtime="00:03:18.09" />
                    <SPLIT distance="250" swimtime="00:04:11.05" />
                    <SPLIT distance="300" swimtime="00:05:04.18" />
                    <SPLIT distance="350" swimtime="00:05:57.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02201" nation="POL" region="01" clubid="2965" name="Uks Shark Rudna">
          <CONTACT name="SZAJNICKI" />
          <ATHLETES>
            <ATHLETE birthdate="1995-07-19" firstname="Katarzyna" gender="F" lastname="Kita" nation="POL" license="102201600048" athleteid="2966">
              <RESULTS>
                <RESULT eventid="1144" points="621" swimtime="00:00:27.80" resultid="7945" heatid="10688" lane="4" entrytime="00:00:27.02" />
                <RESULT eventid="1175" points="443" swimtime="00:02:45.40" resultid="7946" heatid="10717" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:17.66" />
                    <SPLIT distance="150" swimtime="00:02:13.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="421" swimtime="00:00:36.08" resultid="7947" heatid="10739" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1287" points="605" swimtime="00:01:01.54" resultid="7948" heatid="10771" lane="4" entrytime="00:00:59.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="439" swimtime="00:00:32.13" resultid="7949" heatid="10824" lane="3" entrytime="00:00:30.89" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="7950" heatid="10855" lane="3" entrytime="00:02:15.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-02-11" firstname="Agnieszka" gender="F" lastname="Gajdowska" nation="POL" license="102201600071" athleteid="2973">
              <RESULTS>
                <RESULT eventid="1407" points="515" swimtime="00:00:30.46" resultid="9490" heatid="10824" lane="6" entrytime="00:00:31.23" />
                <RESULT eventid="1467" points="498" swimtime="00:02:22.52" resultid="9491" heatid="10855" lane="2" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                    <SPLIT distance="150" swimtime="00:01:45.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="431" swimtime="00:00:39.01" resultid="9492" heatid="10910" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1674" points="470" swimtime="00:05:04.05" resultid="9493" heatid="10934" lane="5" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:12.36" />
                    <SPLIT distance="150" swimtime="00:01:51.76" />
                    <SPLIT distance="200" swimtime="00:02:31.48" />
                    <SPLIT distance="250" swimtime="00:03:10.58" />
                    <SPLIT distance="300" swimtime="00:03:49.96" />
                    <SPLIT distance="350" swimtime="00:04:27.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="571" swimtime="00:00:28.60" resultid="9494" heatid="10688" lane="6" entrytime="00:00:27.98" />
                <RESULT eventid="1175" points="465" swimtime="00:02:42.72" resultid="9495" heatid="10718" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="150" swimtime="00:02:04.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="488" swimtime="00:00:34.35" resultid="9496" heatid="10739" lane="2" entrytime="00:00:33.45" />
                <RESULT eventid="1287" points="584" swimtime="00:01:02.26" resultid="9497" heatid="10771" lane="6" entrytime="00:01:01.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SPCHR" nation="POL" region="MAL" clubid="2835" name="UKS SP 8 Chrzanów">
          <CONTACT city="Chrzanów" email="abalp@poczta.onet.pl" name="Zabrzański  Alfred" phone="692 076 808" state="MAŁ" street="Niepodległości 7 / 46" zip="32 500" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="2842">
              <RESULTS>
                <RESULT eventid="1098" points="173" swimtime="00:13:31.21" resultid="6378" heatid="10670" lane="7" entrytime="00:12:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:01:31.41" />
                    <SPLIT distance="150" swimtime="00:02:20.79" />
                    <SPLIT distance="200" swimtime="00:03:12.86" />
                    <SPLIT distance="250" swimtime="00:04:02.13" />
                    <SPLIT distance="300" swimtime="00:04:52.45" />
                    <SPLIT distance="350" swimtime="00:05:41.06" />
                    <SPLIT distance="400" swimtime="00:06:35.01" />
                    <SPLIT distance="450" swimtime="00:07:26.77" />
                    <SPLIT distance="500" swimtime="00:08:18.51" />
                    <SPLIT distance="550" swimtime="00:09:11.06" />
                    <SPLIT distance="600" swimtime="00:10:02.58" />
                    <SPLIT distance="650" swimtime="00:10:54.41" />
                    <SPLIT distance="700" swimtime="00:11:45.99" />
                    <SPLIT distance="750" swimtime="00:12:39.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="263" swimtime="00:00:32.60" resultid="6379" heatid="10698" lane="4" entrytime="00:00:31.50" entrycourse="SCM" />
                <RESULT eventid="1242" points="182" swimtime="00:00:42.35" resultid="6380" heatid="10744" lane="7" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="1302" points="253" swimtime="00:01:14.13" resultid="6381" heatid="10778" lane="7" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="6382" heatid="10811" lane="2" entrytime="00:01:44.00" entrycourse="SCM" />
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="6383" heatid="10860" lane="0" entrytime="00:02:49.00" entrycourse="SCM" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="6384" heatid="10916" lane="9" entrytime="00:00:44.00" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="6385" heatid="10938" lane="6" entrytime="00:06:21.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02914" nation="POL" region="14" clubid="9083" name="UKS Victoria Józefów">
          <CONTACT email="ali90@o2.pl" name="kowalczyk alicja" />
          <ATHLETES>
            <ATHLETE birthdate="1980-11-08" firstname="Alicja" gender="F" lastname="Kowalczyk-Kędzierska" nation="POL" athleteid="9091">
              <RESULTS>
                <RESULT eventid="1226" points="404" swimtime="00:00:36.59" resultid="9092" heatid="10738" lane="0" entrytime="00:00:38.09" />
                <RESULT eventid="1407" points="367" swimtime="00:00:34.12" resultid="9093" heatid="10823" lane="3" entrytime="00:00:34.09" />
                <RESULT eventid="1437" points="347" swimtime="00:01:22.63" resultid="9094" heatid="10841" lane="3" entrytime="00:01:25.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOKAT" nation="POL" region="SLA" clubid="4122" name="UKS Wodnik 29 Katowice">
          <CONTACT name="Skoczylas" phone="662 297 707" />
          <ATHLETES>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="4123">
              <RESULTS>
                <RESULT eventid="1128" points="294" swimtime="00:21:48.56" resultid="6523" heatid="10678" lane="3" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:17.55" />
                    <SPLIT distance="150" swimtime="00:02:00.31" />
                    <SPLIT distance="200" swimtime="00:02:43.80" />
                    <SPLIT distance="250" swimtime="00:03:27.44" />
                    <SPLIT distance="300" swimtime="00:04:11.08" />
                    <SPLIT distance="350" swimtime="00:04:54.60" />
                    <SPLIT distance="400" swimtime="00:05:38.15" />
                    <SPLIT distance="450" swimtime="00:06:21.65" />
                    <SPLIT distance="500" swimtime="00:07:05.97" />
                    <SPLIT distance="550" swimtime="00:07:50.01" />
                    <SPLIT distance="600" swimtime="00:08:34.02" />
                    <SPLIT distance="650" swimtime="00:09:17.73" />
                    <SPLIT distance="700" swimtime="00:10:02.51" />
                    <SPLIT distance="750" swimtime="00:10:46.17" />
                    <SPLIT distance="800" swimtime="00:11:30.95" />
                    <SPLIT distance="850" swimtime="00:12:15.36" />
                    <SPLIT distance="900" swimtime="00:13:00.01" />
                    <SPLIT distance="950" swimtime="00:13:44.46" />
                    <SPLIT distance="1000" swimtime="00:14:28.86" />
                    <SPLIT distance="1050" swimtime="00:15:13.21" />
                    <SPLIT distance="1100" swimtime="00:15:58.00" />
                    <SPLIT distance="1150" swimtime="00:16:42.27" />
                    <SPLIT distance="1200" swimtime="00:17:26.77" />
                    <SPLIT distance="1250" swimtime="00:18:11.40" />
                    <SPLIT distance="1300" swimtime="00:18:56.39" />
                    <SPLIT distance="1350" swimtime="00:19:41.67" />
                    <SPLIT distance="1400" swimtime="00:20:26.73" />
                    <SPLIT distance="1450" swimtime="00:21:06.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="353" swimtime="00:00:29.57" resultid="6524" heatid="10703" lane="4" entrytime="00:00:28.90" />
                <RESULT eventid="1242" points="274" swimtime="00:00:36.97" resultid="6525" heatid="10747" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1332" points="190" swimtime="00:03:13.92" resultid="6526" heatid="10793" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:28.22" />
                    <SPLIT distance="150" swimtime="00:02:20.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-12-05" firstname="Mariusz" gender="M" lastname="Grelewicz" nation="POL" athleteid="4136">
              <RESULTS>
                <RESULT eventid="1160" points="338" swimtime="00:00:29.99" resultid="6534" heatid="10703" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1638" points="356" swimtime="00:00:37.25" resultid="6535" heatid="10922" lane="6" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-05-18" firstname="Urszula" gender="F" lastname="Walkowicz" nation="POL" athleteid="4143">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat M 85-89 lat" eventid="1144" points="26" swimtime="00:01:19.65" resultid="6539" heatid="10681" lane="1" entrytime="00:01:20.00" />
                <RESULT eventid="1226" status="DNS" swimtime="00:00:00.00" resultid="6540" heatid="10734" lane="7" entrytime="00:01:20.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat mM  85-89  lat" eventid="1287" points="23" swimtime="00:03:01.96" resultid="6541" heatid="10765" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat M  85-89  lat" eventid="1437" points="37" swimtime="00:02:53.11" resultid="6542" heatid="10839" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="30" swimtime="00:06:35.02" resultid="6543" heatid="10893" lane="3" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:36.36" />
                    <SPLIT distance="100" swimtime="00:03:19.97" />
                    <SPLIT distance="150" swimtime="00:05:04.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" status="DNS" swimtime="00:00:00.00" resultid="6544" heatid="10930" lane="5" entrytime="00:13:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="4139">
              <RESULTS>
                <RESULT eventid="1272" points="311" swimtime="00:03:07.41" resultid="6536" heatid="10761" lane="5" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:30.43" />
                    <SPLIT distance="150" swimtime="00:02:19.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="316" swimtime="00:01:23.84" resultid="6537" heatid="10816" lane="1" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="401" swimtime="00:00:35.81" resultid="6538" heatid="10921" lane="4" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-19" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="4128">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="6527" heatid="10697" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1332" status="DNS" swimtime="00:00:00.00" resultid="6529" heatid="10793" lane="0" entrytime="00:03:45.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="6530" heatid="10830" lane="0" entrytime="00:00:34.50" />
                <RESULT eventid="1452" status="DNS" swimtime="00:00:00.00" resultid="6531" heatid="10845" lane="3" entrytime="00:01:35.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="6532" heatid="10886" lane="5" entrytime="00:01:35.00" />
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="6533" heatid="10901" lane="1" entrytime="00:03:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01711" nation="POL" region="11" clubid="3456" name="UKS WODNIK Siemianowice Ślaskie" shortname="UKS WODNIK Siemianowice Ślaski">
          <CONTACT city="Siemianowice Śląskie" email="vivisektor@interia.pl" name="Małyszek Leszek" phone="534033934" state="ŚLĄSK" street="Mikołaja 3" zip="41-106" />
          <ATHLETES>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="3464">
              <RESULTS>
                <RESULT eventid="1128" points="251" swimtime="00:22:59.57" resultid="8044" heatid="10677" lane="7" entrytime="00:22:53.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:24.21" />
                    <SPLIT distance="150" swimtime="00:02:11.13" />
                    <SPLIT distance="200" swimtime="00:02:58.14" />
                    <SPLIT distance="250" swimtime="00:03:43.86" />
                    <SPLIT distance="300" swimtime="00:04:30.35" />
                    <SPLIT distance="350" swimtime="00:05:17.38" />
                    <SPLIT distance="400" swimtime="00:06:03.99" />
                    <SPLIT distance="450" swimtime="00:06:50.83" />
                    <SPLIT distance="500" swimtime="00:07:38.11" />
                    <SPLIT distance="550" swimtime="00:08:23.26" />
                    <SPLIT distance="600" swimtime="00:09:10.16" />
                    <SPLIT distance="650" swimtime="00:09:55.71" />
                    <SPLIT distance="700" swimtime="00:10:39.99" />
                    <SPLIT distance="750" swimtime="00:11:25.73" />
                    <SPLIT distance="800" swimtime="00:12:12.34" />
                    <SPLIT distance="850" swimtime="00:12:58.86" />
                    <SPLIT distance="900" swimtime="00:13:45.12" />
                    <SPLIT distance="950" swimtime="00:14:31.93" />
                    <SPLIT distance="1000" swimtime="00:15:18.55" />
                    <SPLIT distance="1050" swimtime="00:16:04.68" />
                    <SPLIT distance="1100" swimtime="00:16:50.85" />
                    <SPLIT distance="1150" swimtime="00:17:36.34" />
                    <SPLIT distance="1200" swimtime="00:18:21.65" />
                    <SPLIT distance="1250" swimtime="00:19:08.15" />
                    <SPLIT distance="1300" swimtime="00:19:55.07" />
                    <SPLIT distance="1350" swimtime="00:20:41.87" />
                    <SPLIT distance="1400" swimtime="00:21:28.81" />
                    <SPLIT distance="1450" swimtime="00:22:15.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="199" swimtime="00:03:15.12" resultid="8045" heatid="10722" lane="2" entrytime="00:03:10.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                    <SPLIT distance="100" swimtime="00:01:33.74" />
                    <SPLIT distance="150" swimtime="00:02:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="139" swimtime="00:03:35.04" resultid="8046" heatid="10793" lane="1" entrytime="00:03:21.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:42.06" />
                    <SPLIT distance="150" swimtime="00:02:39.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="8047" heatid="10829" lane="1" entrytime="00:00:36.40" />
                <RESULT eventid="1546" status="DNS" swimtime="00:00:00.00" resultid="8048" heatid="10878" lane="5" entrytime="00:06:30.40" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="8049" heatid="10887" lane="1" entrytime="00:01:28.40" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="8050" heatid="10940" lane="1" entrytime="00:05:50.20" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="URWAR" nation="POL" region="14" clubid="4740" name="Ursynów Masters">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1970-01-23" firstname="Michał" gender="M" lastname="Rybarczyk" nation="POL" athleteid="8423">
              <RESULTS>
                <RESULT eventid="1160" points="366" swimtime="00:00:29.21" resultid="8424" heatid="10702" lane="7" entrytime="00:00:29.20" />
                <RESULT eventid="1242" points="124" swimtime="00:00:48.11" resultid="8425" heatid="10744" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1302" points="388" swimtime="00:01:04.31" resultid="8426" heatid="10781" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="318" swimtime="00:00:32.86" resultid="8427" heatid="10830" lane="5" entrytime="00:00:33.84" />
                <RESULT eventid="1482" points="290" swimtime="00:02:34.07" resultid="8428" heatid="10861" lane="8" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="150" swimtime="00:01:56.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="8429" heatid="10887" lane="6" entrytime="00:01:23.00" />
                <RESULT eventid="1695" points="280" swimtime="00:05:36.25" resultid="8430" heatid="10940" lane="6" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:01:18.31" />
                    <SPLIT distance="150" swimtime="00:02:01.57" />
                    <SPLIT distance="200" swimtime="00:02:45.66" />
                    <SPLIT distance="250" swimtime="00:03:30.55" />
                    <SPLIT distance="300" swimtime="00:04:14.39" />
                    <SPLIT distance="350" swimtime="00:04:56.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-03-23" firstname="Ryszard" gender="M" lastname="Rybarczyk" nation="POL" athleteid="4754">
              <RESULTS>
                <RESULT eventid="1160" points="123" swimtime="00:00:42.01" resultid="8431" heatid="10692" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="1242" points="77" swimtime="00:00:56.28" resultid="8432" heatid="10742" lane="9" entrytime="00:00:55.00" />
                <RESULT eventid="1392" points="133" swimtime="00:01:51.74" resultid="8433" heatid="10810" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="55" swimtime="00:02:15.96" resultid="8434" heatid="10844" lane="1" entrytime="00:02:12.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="163" swimtime="00:00:48.30" resultid="8435" heatid="10914" lane="3" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03105" nation="POL" region="05" clubid="4760" name="UTW&quot;Masters&quot; Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1973-03-18" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="503105600018" athleteid="4839">
              <RESULTS>
                <RESULT eventid="1175" points="448" swimtime="00:02:44.71" resultid="8954" heatid="10718" lane="3" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:14.59" />
                    <SPLIT distance="150" swimtime="00:02:03.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="515" swimtime="00:00:33.75" resultid="8955" heatid="10739" lane="3" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1437" points="464" swimtime="00:01:15.02" resultid="8956" heatid="10842" lane="3" entrytime="00:01:13.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="410" swimtime="00:02:46.86" resultid="8957" heatid="10897" lane="3" entrytime="00:02:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                    <SPLIT distance="100" swimtime="00:01:20.41" />
                    <SPLIT distance="150" swimtime="00:02:04.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1922-01-04" firstname="Kazimierz" gender="M" lastname="Mrówczyński" nation="POL" license="503105700021" athleteid="8880">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Europy Masters Mężczyzn w  kat O 95-99 lat" eventid="1160" points="34" swimtime="00:01:04.37" resultid="8881" heatid="10690" lane="4" entrytime="00:01:01.00" entrycourse="LCM" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="8882" heatid="10773" lane="8" entrytime="00:02:40.00" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Europy Masters  Mężczyzn w  kat O  95-99  lat, międzyczas na 100 m dow lepszy od Rekordu Europy Masters w kat. O 95-99 lat" eventid="1482" points="27" swimtime="00:05:36.99" resultid="8883" heatid="10856" lane="3" entrytime="00:05:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.40" />
                    <SPLIT distance="100" swimtime="00:02:41.94" />
                    <SPLIT distance="150" swimtime="00:04:12.03" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Europy, nieoficjalny Rekord Polski" eventid="1638" points="38" swimtime="00:01:18.50" resultid="8884" heatid="10913" lane="9" entrytime="00:01:18.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105700034" athleteid="4828">
              <RESULTS>
                <RESULT eventid="1098" points="113" swimtime="00:15:32.90" resultid="8945" heatid="10669" lane="6" entrytime="00:17:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.40" />
                    <SPLIT distance="100" swimtime="00:01:46.73" />
                    <SPLIT distance="150" swimtime="00:02:46.13" />
                    <SPLIT distance="200" swimtime="00:03:45.59" />
                    <SPLIT distance="250" swimtime="00:04:42.95" />
                    <SPLIT distance="300" swimtime="00:05:41.62" />
                    <SPLIT distance="350" swimtime="00:06:40.78" />
                    <SPLIT distance="400" swimtime="00:07:38.68" />
                    <SPLIT distance="450" swimtime="00:08:38.24" />
                    <SPLIT distance="500" swimtime="00:09:38.35" />
                    <SPLIT distance="550" swimtime="00:10:38.30" />
                    <SPLIT distance="600" swimtime="00:11:38.10" />
                    <SPLIT distance="650" swimtime="00:12:38.41" />
                    <SPLIT distance="700" swimtime="00:13:38.53" />
                    <SPLIT distance="750" swimtime="00:14:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="199" swimtime="00:03:37.29" resultid="8946" heatid="10757" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.51" />
                    <SPLIT distance="100" swimtime="00:01:46.32" />
                    <SPLIT distance="150" swimtime="00:02:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="200" swimtime="00:01:37.58" resultid="8947" heatid="10809" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="263" swimtime="00:00:41.23" resultid="8948" heatid="10916" lane="3" entrytime="00:00:42.30" entrycourse="LCM" />
                <RESULT eventid="1695" points="110" swimtime="00:07:39.18" resultid="8949" heatid="10936" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.92" />
                    <SPLIT distance="100" swimtime="00:01:45.27" />
                    <SPLIT distance="150" swimtime="00:02:45.41" />
                    <SPLIT distance="200" swimtime="00:03:45.83" />
                    <SPLIT distance="250" swimtime="00:04:45.64" />
                    <SPLIT distance="300" swimtime="00:05:46.83" />
                    <SPLIT distance="350" swimtime="00:06:46.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="Błasiak" nation="POL" license="503105700050" athleteid="8894">
              <RESULTS>
                <RESULT eventid="1160" points="137" swimtime="00:00:40.47" resultid="8895" heatid="10692" lane="4" entrytime="00:00:39.42" entrycourse="LCM" />
                <RESULT eventid="1190" points="79" swimtime="00:04:24.70" resultid="8896" heatid="10720" lane="0" entrytime="00:04:27.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.71" />
                    <SPLIT distance="100" swimtime="00:02:09.98" />
                    <SPLIT distance="150" swimtime="00:03:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="122" swimtime="00:01:34.36" resultid="8897" heatid="10774" lane="0" entrytime="00:01:35.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="51" swimtime="00:05:00.13" resultid="8898" heatid="10792" lane="9" entrytime="00:04:56.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.91" />
                    <SPLIT distance="100" swimtime="00:02:24.73" />
                    <SPLIT distance="150" swimtime="00:03:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="94" swimtime="00:03:43.80" resultid="8899" heatid="10857" lane="2" entrytime="00:03:35.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="80" swimtime="00:09:23.85" resultid="8900" heatid="10876" lane="4" entrytime="00:09:10.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.22" />
                    <SPLIT distance="100" swimtime="00:02:28.02" />
                    <SPLIT distance="150" swimtime="00:03:41.57" />
                    <SPLIT distance="200" swimtime="00:04:53.62" />
                    <SPLIT distance="250" swimtime="00:06:14.32" />
                    <SPLIT distance="300" swimtime="00:07:30.76" />
                    <SPLIT distance="350" swimtime="00:08:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="39" swimtime="00:02:26.90" resultid="8901" heatid="10885" lane="3" entrytime="00:02:14.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="97" swimtime="00:07:57.36" resultid="8902" heatid="10936" lane="3" entrytime="00:07:51.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.49" />
                    <SPLIT distance="100" swimtime="00:01:51.13" />
                    <SPLIT distance="150" swimtime="00:02:54.14" />
                    <SPLIT distance="200" swimtime="00:03:56.63" />
                    <SPLIT distance="250" swimtime="00:05:00.60" />
                    <SPLIT distance="300" swimtime="00:06:02.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-27" firstname="Natalia" gender="F" lastname="Szczęsnowicz" nation="POL" license="503105600052" athleteid="8912">
              <RESULTS>
                <RESULT eventid="1144" points="385" swimtime="00:00:32.60" resultid="8913" heatid="10687" lane="5" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1226" status="DNS" swimtime="00:00:00.00" resultid="8914" heatid="10734" lane="8" />
                <RESULT eventid="1376" points="366" swimtime="00:01:29.89" resultid="8915" heatid="10803" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="338" swimtime="00:00:35.07" resultid="8916" heatid="10823" lane="7" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1623" points="394" swimtime="00:00:40.21" resultid="8917" heatid="10911" lane="9" entrytime="00:00:38.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-05-25" firstname="Włodzimierz" gender="M" lastname="Łatecki" nation="POL" license="503105700032" athleteid="8885">
              <RESULTS>
                <RESULT eventid="1190" points="55" swimtime="00:04:59.47" resultid="8886" heatid="10719" lane="3" entrytime="00:05:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.78" />
                    <SPLIT distance="100" swimtime="00:02:32.19" />
                    <SPLIT distance="150" swimtime="00:03:59.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="41" swimtime="00:05:20.84" resultid="8887" heatid="10791" lane="4" entrytime="00:05:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.44" />
                    <SPLIT distance="100" swimtime="00:02:32.91" />
                    <SPLIT distance="150" swimtime="00:03:58.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="57" swimtime="00:10:32.00" resultid="8888" heatid="10876" lane="5" entrytime="00:09:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.82" />
                    <SPLIT distance="100" swimtime="00:02:32.95" />
                    <SPLIT distance="150" swimtime="00:03:59.21" />
                    <SPLIT distance="200" swimtime="00:05:30.63" />
                    <SPLIT distance="250" swimtime="00:06:56.83" />
                    <SPLIT distance="300" swimtime="00:08:26.81" />
                    <SPLIT distance="350" swimtime="00:09:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="76" swimtime="00:08:39.24" resultid="8889" heatid="10936" lane="2" entrytime="00:08:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.77" />
                    <SPLIT distance="100" swimtime="00:01:56.78" />
                    <SPLIT distance="150" swimtime="00:03:05.11" />
                    <SPLIT distance="200" swimtime="00:04:12.26" />
                    <SPLIT distance="250" swimtime="00:05:21.23" />
                    <SPLIT distance="300" swimtime="00:06:29.30" />
                    <SPLIT distance="350" swimtime="00:07:36.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-02-07" firstname="Krzysztof" gender="M" lastname="Wojciechowski" nation="POL" license="503105700024" athleteid="4771">
              <RESULTS>
                <RESULT eventid="1190" points="151" swimtime="00:03:33.90" resultid="8890" heatid="10721" lane="9" entrytime="00:03:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                    <SPLIT distance="100" swimtime="00:01:46.80" />
                    <SPLIT distance="150" swimtime="00:02:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="195" swimtime="00:03:38.92" resultid="8891" heatid="10759" lane="7" entrytime="00:03:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                    <SPLIT distance="100" swimtime="00:01:45.72" />
                    <SPLIT distance="150" swimtime="00:02:44.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="214" swimtime="00:01:35.49" resultid="8892" heatid="10813" lane="8" entrytime="00:01:34.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="275" swimtime="00:00:40.60" resultid="8893" heatid="10917" lane="2" entrytime="00:00:41.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105700026" athleteid="4804">
              <RESULTS>
                <RESULT eventid="1160" points="254" swimtime="00:00:32.98" resultid="8922" heatid="10696" lane="5" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1302" points="232" swimtime="00:01:16.28" resultid="8923" heatid="10776" lane="4" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" status="DNS" swimtime="00:00:00.00" resultid="8924" heatid="10791" lane="2" />
                <RESULT eventid="1422" points="217" swimtime="00:00:37.29" resultid="8925" heatid="10829" lane="9" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="1546" points="99" swimtime="00:08:46.62" resultid="8926" heatid="10876" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.47" />
                    <SPLIT distance="100" swimtime="00:02:18.23" />
                    <SPLIT distance="150" swimtime="00:03:30.46" />
                    <SPLIT distance="200" swimtime="00:04:38.72" />
                    <SPLIT distance="250" swimtime="00:05:55.71" />
                    <SPLIT distance="300" swimtime="00:07:11.83" />
                    <SPLIT distance="350" swimtime="00:08:01.71" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1578" points="131" swimtime="00:01:37.97" resultid="8927" heatid="10886" lane="6" entrytime="00:01:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="503105700038" athleteid="8918">
              <RESULTS>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="8919" heatid="10758" lane="3" entrytime="00:03:47.00" entrycourse="LCM" />
                <RESULT eventid="1392" points="206" swimtime="00:01:36.73" resultid="8920" heatid="10812" lane="5" entrytime="00:01:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="265" swimtime="00:00:41.11" resultid="8921" heatid="10916" lane="6" entrytime="00:00:42.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105600028" athleteid="8958">
              <RESULTS>
                <RESULT eventid="1175" points="416" swimtime="00:02:48.89" resultid="8959" heatid="10717" lane="3" entrytime="00:02:47.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:18.27" />
                    <SPLIT distance="150" swimtime="00:02:08.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="342" swimtime="00:00:38.67" resultid="8960" heatid="10739" lane="8" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1317" points="308" swimtime="00:03:00.23" resultid="8961" heatid="10790" lane="2" entrytime="00:03:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:01:26.24" />
                    <SPLIT distance="150" swimtime="00:02:12.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="423" swimtime="00:00:32.52" resultid="8962" heatid="10823" lane="5" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1437" points="332" swimtime="00:01:23.93" resultid="8963" heatid="10842" lane="2" entrytime="00:01:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="433" swimtime="00:01:13.30" resultid="8964" heatid="10883" lane="2" entrytime="00:01:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" status="DNS" swimtime="00:00:00.00" resultid="8965" heatid="10897" lane="8" entrytime="00:02:50.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-16" firstname="Adrian" gender="M" lastname="Styrzyński" nation="POL" license="503105700033" athleteid="8966">
              <RESULTS>
                <RESULT eventid="1160" points="565" swimtime="00:00:25.29" resultid="8967" heatid="10711" lane="3" entrytime="00:00:24.20" entrycourse="LCM" />
                <RESULT eventid="1302" points="577" swimtime="00:00:56.33" resultid="8968" heatid="10788" lane="1" entrytime="00:00:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="495" swimtime="00:01:12.20" resultid="8969" heatid="10819" lane="3" entrytime="00:01:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="8970" heatid="10866" lane="3" entrytime="00:01:59.99" entrycourse="LCM" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="8971" heatid="10892" lane="6" entrytime="00:00:59.00" entrycourse="LCM" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="8972" heatid="10926" lane="3" entrytime="00:00:29.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-01" firstname="Waldemar" gender="M" lastname="Jagiełło" nation="POL" license="503105700036" athleteid="8903">
              <RESULTS>
                <RESULT eventid="1160" points="498" swimtime="00:00:26.37" resultid="8904" heatid="10705" lane="4" entrytime="00:00:27.65" entrycourse="LCM" />
                <RESULT eventid="1190" points="397" swimtime="00:02:34.99" resultid="8905" heatid="10728" lane="8" entrytime="00:02:36.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:02:00.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="431" swimtime="00:02:48.07" resultid="8906" heatid="10763" lane="5" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:16.34" />
                    <SPLIT distance="150" swimtime="00:02:01.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="492" swimtime="00:00:59.41" resultid="8907" heatid="10785" lane="3" entrytime="00:00:59.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="447" swimtime="00:01:14.68" resultid="8908" heatid="10818" lane="7" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="457" swimtime="00:00:29.11" resultid="8909" heatid="10835" lane="1" entrytime="00:00:29.65" entrycourse="LCM" />
                <RESULT eventid="1578" points="399" swimtime="00:01:07.67" resultid="8910" heatid="10890" lane="1" entrytime="00:01:09.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="533" swimtime="00:00:32.58" resultid="8911" heatid="10925" lane="1" entrytime="00:00:32.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="Ewa" gender="F" lastname="Stępień" nation="POL" license="503105600029" athleteid="8936">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat G 55-59 lat" eventid="1144" points="399" swimtime="00:00:32.21" resultid="8937" heatid="10685" lane="2" entrytime="00:00:34.02" entrycourse="LCM" />
                <RESULT eventid="1175" points="320" swimtime="00:03:04.38" resultid="8938" heatid="10716" lane="5" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                    <SPLIT distance="100" swimtime="00:01:27.65" />
                    <SPLIT distance="150" swimtime="00:02:19.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="316" swimtime="00:03:24.19" resultid="8939" heatid="10755" lane="2" entrytime="00:03:20.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                    <SPLIT distance="100" swimtime="00:01:36.34" />
                    <SPLIT distance="150" swimtime="00:02:29.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat G  55-59  lat" eventid="1287" points="333" swimtime="00:01:15.07" resultid="8940" heatid="10770" lane="0" entrytime="00:01:14.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat G  55-59  lat" eventid="1376" points="371" swimtime="00:01:29.50" resultid="8941" heatid="10807" lane="5" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="278" swimtime="00:02:52.93" resultid="8942" heatid="10854" lane="0" entrytime="00:02:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:01:21.35" />
                    <SPLIT distance="150" swimtime="00:02:06.88" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1623" points="380" swimtime="00:00:40.69" resultid="8943" heatid="10910" lane="8" entrytime="00:00:40.30" entrycourse="LCM" />
                <RESULT eventid="1674" status="DNS" swimtime="00:00:00.00" resultid="8944" heatid="10933" lane="3" entrytime="00:05:55.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-25" firstname="Michał" gender="M" lastname="Woźniak" nation="POL" license="503105700039" athleteid="8973">
              <RESULTS>
                <RESULT eventid="1098" points="337" swimtime="00:10:49.18" resultid="8974" heatid="10673" lane="3" entrytime="00:09:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:51.47" />
                    <SPLIT distance="200" swimtime="00:02:31.89" />
                    <SPLIT distance="250" swimtime="00:03:12.65" />
                    <SPLIT distance="300" swimtime="00:03:53.14" />
                    <SPLIT distance="350" swimtime="00:04:34.72" />
                    <SPLIT distance="400" swimtime="00:05:16.38" />
                    <SPLIT distance="450" swimtime="00:05:58.22" />
                    <SPLIT distance="500" swimtime="00:06:39.70" />
                    <SPLIT distance="550" swimtime="00:07:21.41" />
                    <SPLIT distance="600" swimtime="00:08:02.87" />
                    <SPLIT distance="650" swimtime="00:08:44.89" />
                    <SPLIT distance="700" swimtime="00:09:26.34" />
                    <SPLIT distance="750" swimtime="00:10:08.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="8975" heatid="10709" lane="3" entrytime="00:00:26.00" entrycourse="LCM" />
                <RESULT eventid="1242" points="427" swimtime="00:00:31.90" resultid="8976" heatid="10751" lane="9" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1452" points="432" swimtime="00:01:08.54" resultid="8977" heatid="10849" lane="5" entrytime="00:01:07.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="394" swimtime="00:02:32.61" resultid="8978" heatid="10904" lane="6" entrytime="00:02:26.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:13.34" />
                    <SPLIT distance="150" swimtime="00:01:53.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-23" firstname="Tomasz" gender="M" lastname="Cajdler" nation="POL" license="503105700035" athleteid="4834">
              <RESULTS>
                <RESULT eventid="1160" points="250" swimtime="00:00:33.19" resultid="8950" heatid="10697" lane="8" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1302" points="231" swimtime="00:01:16.39" resultid="8951" heatid="10776" lane="5" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="171" swimtime="00:01:42.88" resultid="8952" heatid="10812" lane="6" entrytime="00:01:36.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="227" swimtime="00:00:43.25" resultid="8953" heatid="10916" lane="1" entrytime="00:00:43.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105600030" athleteid="8928">
              <RESULTS>
                <RESULT eventid="1144" points="343" swimtime="00:00:33.87" resultid="8929" heatid="10685" lane="3" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat G  55-59  lat" eventid="1226" points="317" swimtime="00:00:39.65" resultid="8930" heatid="10738" lane="9" entrytime="00:00:38.30" entrycourse="LCM" />
                <RESULT eventid="1317" points="196" swimtime="00:03:29.64" resultid="8931" heatid="10790" lane="7" entrytime="00:03:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:41.17" />
                    <SPLIT distance="150" swimtime="00:02:35.63" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat G  55-59  lat" eventid="1407" points="330" swimtime="00:00:35.32" resultid="8932" heatid="10823" lane="9" entrytime="00:00:36.20" entrycourse="LCM" />
                <RESULT eventid="1437" points="245" swimtime="00:01:32.77" resultid="8933" heatid="10841" lane="6" entrytime="00:01:26.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1562" points="249" swimtime="00:01:28.10" resultid="8934" heatid="10884" lane="9" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="212" swimtime="00:06:36.45" resultid="8935" heatid="10933" lane="4" entrytime="00:05:54.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:29.25" />
                    <SPLIT distance="150" swimtime="00:02:19.64" />
                    <SPLIT distance="200" swimtime="00:03:13.21" />
                    <SPLIT distance="250" swimtime="00:04:05.15" />
                    <SPLIT distance="300" swimtime="00:04:56.00" />
                    <SPLIT distance="350" swimtime="00:05:48.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105700027" athleteid="8979">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Mężczyzn w  kat H 60-64 lata" eventid="1098" points="256" swimtime="00:11:51.76" resultid="8980" heatid="10671" lane="0" entrytime="00:11:58.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:02:01.42" />
                    <SPLIT distance="200" swimtime="00:02:45.41" />
                    <SPLIT distance="250" swimtime="00:03:30.72" />
                    <SPLIT distance="300" swimtime="00:04:15.83" />
                    <SPLIT distance="350" swimtime="00:05:01.18" />
                    <SPLIT distance="400" swimtime="00:05:46.95" />
                    <SPLIT distance="450" swimtime="00:06:32.87" />
                    <SPLIT distance="500" swimtime="00:07:19.45" />
                    <SPLIT distance="550" swimtime="00:08:05.40" />
                    <SPLIT distance="600" swimtime="00:08:52.28" />
                    <SPLIT distance="650" swimtime="00:09:39.69" />
                    <SPLIT distance="700" swimtime="00:10:25.29" />
                    <SPLIT distance="750" swimtime="00:11:09.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="307" swimtime="00:00:30.97" resultid="8981" heatid="10699" lane="8" entrytime="00:00:31.00" entrycourse="LCM" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="8982" heatid="10723" lane="3" entrytime="00:03:00.00" entrycourse="LCM" />
                <RESULT eventid="1242" points="289" swimtime="00:00:36.36" resultid="8983" heatid="10746" lane="5" entrytime="00:00:36.30" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn w  kat H  60-64  lata" eventid="1332" points="215" swimtime="00:03:06.09" resultid="8984" heatid="10793" lane="5" entrytime="00:03:12.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                    <SPLIT distance="100" swimtime="00:01:30.08" />
                    <SPLIT distance="150" swimtime="00:02:18.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="334" swimtime="00:00:32.31" resultid="8985" heatid="10832" lane="8" entrytime="00:00:32.28" entrycourse="LCM" />
                <RESULT eventid="1546" points="234" swimtime="00:06:35.51" resultid="8986" heatid="10879" lane="9" entrytime="00:06:27.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                    <SPLIT distance="100" swimtime="00:01:33.89" />
                    <SPLIT distance="150" swimtime="00:02:25.47" />
                    <SPLIT distance="200" swimtime="00:03:16.21" />
                    <SPLIT distance="250" swimtime="00:04:17.63" />
                    <SPLIT distance="300" swimtime="00:05:17.60" />
                    <SPLIT distance="350" swimtime="00:05:57.78" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1578" points="257" swimtime="00:01:18.32" resultid="8987" heatid="10887" lane="4" entrytime="00:01:21.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1695" points="276" swimtime="00:05:37.98" resultid="8988" heatid="10941" lane="1" entrytime="00:05:39.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                    <SPLIT distance="200" swimtime="00:02:44.78" />
                    <SPLIT distance="250" swimtime="00:03:29.74" />
                    <SPLIT distance="300" swimtime="00:04:13.68" />
                    <SPLIT distance="350" swimtime="00:04:57.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-03" firstname="Stanisław" gender="M" lastname="Sikorski" nation="POL" license="503105700054" athleteid="8989">
              <RESULTS>
                <RESULT eventid="1242" points="94" swimtime="00:00:52.85" resultid="8990" heatid="10742" lane="3" entrytime="00:00:50.00" entrycourse="LCM" />
                <RESULT eventid="1392" points="117" swimtime="00:01:56.76" resultid="8991" heatid="10810" lane="9" entrytime="00:02:04.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="57" swimtime="00:02:14.72" resultid="8992" heatid="10844" lane="6" entrytime="00:02:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="155" swimtime="00:00:49.14" resultid="8993" heatid="10914" lane="2" entrytime="00:00:50.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="450" swimtime="00:02:01.90" resultid="8995" heatid="10802" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:04.60" />
                    <SPLIT distance="150" swimtime="00:01:30.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8973" number="1" />
                    <RELAYPOSITION athleteid="8903" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="8966" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="8979" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" points="455" swimtime="00:01:50.29" resultid="8996" heatid="10872" lane="8" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                    <SPLIT distance="100" swimtime="00:00:53.99" />
                    <SPLIT distance="150" swimtime="00:01:25.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8903" number="1" />
                    <RELAYPOSITION athleteid="8973" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="8979" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="8966" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1368" points="188" swimtime="00:02:43.04" resultid="8997" heatid="10800" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.97" />
                    <SPLIT distance="100" swimtime="00:01:27.49" />
                    <SPLIT distance="150" swimtime="00:02:09.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4771" number="1" />
                    <RELAYPOSITION athleteid="4828" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4804" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4834" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1518" points="222" swimtime="00:02:20.06" resultid="8998" heatid="10870" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:11.02" />
                    <SPLIT distance="150" swimtime="00:01:46.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4804" number="1" />
                    <RELAYPOSITION athleteid="4828" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4771" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4834" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  w  kat D  200-239  lata" eventid="1347" points="413" swimtime="00:02:22.68" resultid="8999" heatid="10798" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:15.14" />
                    <SPLIT distance="150" swimtime="00:01:49.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4839" number="1" />
                    <RELAYPOSITION athleteid="8936" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="8928" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="8958" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1497" points="419" swimtime="00:02:08.93" resultid="9000" heatid="10868" lane="9" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="100" swimtime="00:01:07.13" />
                    <SPLIT distance="150" swimtime="00:01:38.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8936" number="1" />
                    <RELAYPOSITION athleteid="8928" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="8958" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4839" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:26.50" resultid="8994" heatid="10928" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                    <SPLIT distance="100" swimtime="00:01:20.42" />
                    <SPLIT distance="150" swimtime="00:01:52.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8928" number="1" />
                    <RELAYPOSITION athleteid="8936" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="8979" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4804" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:01:57.50" resultid="9002" heatid="10733" lane="0" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                    <SPLIT distance="100" swimtime="00:01:03.13" />
                    <SPLIT distance="150" swimtime="00:01:29.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8958" number="1" />
                    <RELAYPOSITION athleteid="8973" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4839" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="8903" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1653" swimtime="00:02:07.39" resultid="9001" heatid="10929" lane="5" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:04.89" />
                    <SPLIT distance="150" swimtime="00:01:37.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8973" number="1" />
                    <RELAYPOSITION athleteid="8903" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="8958" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4839" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:11.11" resultid="9003" heatid="10732" lane="7" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:07.96" />
                    <SPLIT distance="150" swimtime="00:01:40.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4804" number="1" />
                    <RELAYPOSITION athleteid="8928" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="8936" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="8979" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="USOST" nation="POL" region="14" clubid="6069" name="Uśks Ostrołęka">
          <CONTACT name="UŚKS OSTROŁĘKA" />
          <ATHLETES>
            <ATHLETE birthdate="1990-12-06" firstname="Adam" gender="M" lastname="Janczewski" nation="POL" license="501914700035" athleteid="6070">
              <RESULTS>
                <RESULT eventid="1098" points="333" swimtime="00:10:51.94" resultid="7767" heatid="10672" lane="3" entrytime="00:10:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:13.94" />
                    <SPLIT distance="150" swimtime="00:01:53.84" />
                    <SPLIT distance="200" swimtime="00:02:34.14" />
                    <SPLIT distance="250" swimtime="00:03:14.31" />
                    <SPLIT distance="300" swimtime="00:03:55.24" />
                    <SPLIT distance="350" swimtime="00:04:36.03" />
                    <SPLIT distance="400" swimtime="00:05:16.93" />
                    <SPLIT distance="450" swimtime="00:05:58.24" />
                    <SPLIT distance="500" swimtime="00:06:40.14" />
                    <SPLIT distance="550" swimtime="00:07:22.50" />
                    <SPLIT distance="600" swimtime="00:08:04.68" />
                    <SPLIT distance="650" swimtime="00:08:47.09" />
                    <SPLIT distance="700" swimtime="00:09:29.57" />
                    <SPLIT distance="750" swimtime="00:10:11.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="445" swimtime="00:02:29.22" resultid="7768" heatid="10729" lane="4" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                    <SPLIT distance="100" swimtime="00:01:10.81" />
                    <SPLIT distance="150" swimtime="00:01:56.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="7769" heatid="10944" lane="0" entrytime="00:04:59.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAELB" nation="POL" region="WAR" clubid="4066" name="Victory Masters Elbląg">
          <CONTACT city="Elbląg" name="Latecki Grzegorz" street="Łokietka" street2="45" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner-Mateusiak" nation="POL" athleteid="4098">
              <RESULTS>
                <RESULT eventid="1059" points="54" swimtime="00:21:20.67" resultid="6454" heatid="10666" lane="1" entrytime="00:17:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.84" />
                    <SPLIT distance="100" swimtime="00:02:23.85" />
                    <SPLIT distance="150" swimtime="00:03:45.44" />
                    <SPLIT distance="200" swimtime="00:05:09.06" />
                    <SPLIT distance="250" swimtime="00:06:29.52" />
                    <SPLIT distance="300" swimtime="00:07:51.80" />
                    <SPLIT distance="350" swimtime="00:09:10.82" />
                    <SPLIT distance="400" swimtime="00:10:32.09" />
                    <SPLIT distance="450" swimtime="00:11:37.00" />
                    <SPLIT distance="550" swimtime="00:11:53.16" />
                    <SPLIT distance="600" swimtime="00:13:15.81" />
                    <SPLIT distance="650" swimtime="00:14:36.49" />
                    <SPLIT distance="700" swimtime="00:15:59.31" />
                    <SPLIT distance="750" swimtime="00:17:18.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1226" points="63" swimtime="00:01:07.70" resultid="6455" heatid="10734" lane="2" entrytime="00:01:06.77" />
                <RESULT comment="O 4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1257" status="DSQ" swimtime="00:05:48.33" resultid="6456" heatid="10752" lane="5" entrytime="00:05:35.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.82" />
                    <SPLIT distance="100" swimtime="00:02:51.42" />
                    <SPLIT distance="150" swimtime="00:04:18.71" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 14 - Praca nóg  w płaszczyźnie pionowej w dół /z wyjątkiem jednego ruchu po starcie i nawrocie/" eventid="1376" status="DSQ" swimtime="00:02:48.05" resultid="6457" heatid="10803" lane="2" entrytime="00:02:42.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="53" swimtime="00:02:34.72" resultid="6458" heatid="10839" lane="7" entrytime="00:02:28.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="56" swimtime="00:05:23.01" resultid="6459" heatid="10893" lane="4" entrytime="00:05:27.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.68" />
                    <SPLIT distance="100" swimtime="00:02:41.29" />
                    <SPLIT distance="150" swimtime="00:04:03.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="56" swimtime="00:10:16.94" resultid="6460" heatid="10931" lane="0" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.58" />
                    <SPLIT distance="100" swimtime="00:02:24.11" />
                    <SPLIT distance="150" swimtime="00:03:43.25" />
                    <SPLIT distance="200" swimtime="00:05:01.44" />
                    <SPLIT distance="250" swimtime="00:06:17.83" />
                    <SPLIT distance="300" swimtime="00:07:37.27" />
                    <SPLIT distance="350" swimtime="00:08:57.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="Karaś" nation="POL" athleteid="4090">
              <RESULTS>
                <RESULT eventid="1059" points="154" swimtime="00:15:04.09" resultid="6447" heatid="10667" lane="9" entrytime="00:14:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.72" />
                    <SPLIT distance="100" swimtime="00:01:46.60" />
                    <SPLIT distance="150" swimtime="00:02:42.88" />
                    <SPLIT distance="200" swimtime="00:03:39.34" />
                    <SPLIT distance="250" swimtime="00:04:36.49" />
                    <SPLIT distance="300" swimtime="00:05:33.41" />
                    <SPLIT distance="350" swimtime="00:06:30.64" />
                    <SPLIT distance="400" swimtime="00:07:28.11" />
                    <SPLIT distance="450" swimtime="00:08:25.70" />
                    <SPLIT distance="500" swimtime="00:09:23.19" />
                    <SPLIT distance="550" swimtime="00:10:21.54" />
                    <SPLIT distance="600" swimtime="00:11:20.00" />
                    <SPLIT distance="650" swimtime="00:12:16.99" />
                    <SPLIT distance="700" swimtime="00:13:15.24" />
                    <SPLIT distance="750" swimtime="00:14:10.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="112" swimtime="00:04:21.46" resultid="6448" heatid="10713" lane="1" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.07" />
                    <SPLIT distance="100" swimtime="00:02:06.18" />
                    <SPLIT distance="150" swimtime="00:03:26.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1317" points="103" swimtime="00:04:19.74" resultid="6449" heatid="10789" lane="4" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.12" />
                    <SPLIT distance="100" swimtime="00:02:03.63" />
                    <SPLIT distance="150" swimtime="00:03:12.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="151" swimtime="00:03:32.01" resultid="6450" heatid="10852" lane="8" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                    <SPLIT distance="100" swimtime="00:01:42.47" />
                    <SPLIT distance="150" swimtime="00:02:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 14 - Praca nóg  w płaszczyźnie pionowej w dół /z wyjątkiem jednego ruchu po starcie i nawrocie/" eventid="1525" status="DSQ" swimtime="00:08:50.42" resultid="6451" heatid="10873" lane="5" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.93" />
                    <SPLIT distance="100" swimtime="00:02:02.72" />
                    <SPLIT distance="150" swimtime="00:03:11.67" />
                    <SPLIT distance="200" swimtime="00:04:21.67" />
                    <SPLIT distance="250" swimtime="00:05:42.02" />
                    <SPLIT distance="300" swimtime="00:07:01.92" />
                    <SPLIT distance="350" swimtime="00:07:57.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="97" swimtime="00:02:00.70" resultid="6452" heatid="10883" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="155" swimtime="00:07:19.88" resultid="6453" heatid="10932" lane="9" entrytime="00:07:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.85" />
                    <SPLIT distance="100" swimtime="00:01:45.97" />
                    <SPLIT distance="150" swimtime="00:02:41.87" />
                    <SPLIT distance="200" swimtime="00:03:38.15" />
                    <SPLIT distance="250" swimtime="00:04:34.67" />
                    <SPLIT distance="300" swimtime="00:05:30.63" />
                    <SPLIT distance="350" swimtime="00:06:26.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-12" firstname="Grzegorz" gender="M" lastname="Latecki" nation="POL" athleteid="4075">
              <RESULTS>
                <RESULT eventid="1160" points="408" swimtime="00:00:28.18" resultid="6434" heatid="10704" lane="8" entrytime="00:00:28.70" />
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="6436" heatid="10748" lane="2" entrytime="00:00:33.60" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="6437" heatid="10783" lane="3" entrytime="00:01:02.90" />
                <RESULT eventid="1422" points="445" swimtime="00:00:29.36" resultid="6438" heatid="10834" lane="1" entrytime="00:00:30.30" />
                <RESULT eventid="1546" points="328" swimtime="00:05:53.40" resultid="6439" heatid="10879" lane="3" entrytime="00:06:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                    <SPLIT distance="150" swimtime="00:02:05.08" />
                    <SPLIT distance="200" swimtime="00:02:51.70" />
                    <SPLIT distance="250" swimtime="00:03:42.64" />
                    <SPLIT distance="300" swimtime="00:04:35.37" />
                    <SPLIT distance="350" swimtime="00:05:14.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="371" swimtime="00:01:09.28" resultid="6440" heatid="10889" lane="3" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="6441" heatid="10920" lane="5" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="4084">
              <RESULTS>
                <RESULT eventid="1059" points="143" swimtime="00:15:27.05" resultid="6442" heatid="10667" lane="8" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.97" />
                    <SPLIT distance="100" swimtime="00:01:51.35" />
                    <SPLIT distance="150" swimtime="00:02:50.45" />
                    <SPLIT distance="200" swimtime="00:03:49.87" />
                    <SPLIT distance="250" swimtime="00:04:49.61" />
                    <SPLIT distance="300" swimtime="00:05:49.27" />
                    <SPLIT distance="350" swimtime="00:06:48.10" />
                    <SPLIT distance="400" swimtime="00:07:47.56" />
                    <SPLIT distance="450" swimtime="00:08:46.11" />
                    <SPLIT distance="500" swimtime="00:09:44.55" />
                    <SPLIT distance="550" swimtime="00:10:42.57" />
                    <SPLIT distance="600" swimtime="00:11:39.80" />
                    <SPLIT distance="650" swimtime="00:12:37.03" />
                    <SPLIT distance="700" swimtime="00:13:34.88" />
                    <SPLIT distance="750" swimtime="00:14:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="149" swimtime="00:00:44.70" resultid="6443" heatid="10682" lane="1" entrytime="00:00:43.72" />
                <RESULT eventid="1287" points="141" swimtime="00:01:39.87" resultid="6444" heatid="10766" lane="3" entrytime="00:01:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="146" swimtime="00:03:34.49" resultid="6445" heatid="10852" lane="9" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.51" />
                    <SPLIT distance="100" swimtime="00:01:45.54" />
                    <SPLIT distance="150" swimtime="00:02:42.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="143" swimtime="00:07:32.01" resultid="6446" heatid="10932" lane="8" entrytime="00:07:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.76" />
                    <SPLIT distance="100" swimtime="00:01:50.30" />
                    <SPLIT distance="150" swimtime="00:02:49.32" />
                    <SPLIT distance="200" swimtime="00:03:48.40" />
                    <SPLIT distance="250" swimtime="00:04:46.73" />
                    <SPLIT distance="300" swimtime="00:05:44.08" />
                    <SPLIT distance="350" swimtime="00:06:41.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-06" firstname="Andrzej" gender="M" lastname="Pasieczny" nation="POL" athleteid="4067">
              <RESULTS>
                <RESULT eventid="1160" points="379" swimtime="00:00:28.87" resultid="6427" heatid="10704" lane="0" entrytime="00:00:28.72" />
                <RESULT eventid="1190" points="423" swimtime="00:02:31.80" resultid="6428" heatid="10728" lane="9" entrytime="00:02:37.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="150" swimtime="00:01:57.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="424" swimtime="00:01:02.41" resultid="6429" heatid="10783" lane="9" entrytime="00:01:03.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="400" swimtime="00:00:30.43" resultid="6430" heatid="10833" lane="5" entrytime="00:00:30.56" />
                <RESULT eventid="1482" points="432" swimtime="00:02:14.83" resultid="6431" heatid="10865" lane="9" entrytime="00:02:14.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:05.40" />
                    <SPLIT distance="150" swimtime="00:01:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="425" swimtime="00:01:06.25" resultid="6432" heatid="10890" lane="5" entrytime="00:01:05.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1695" points="442" swimtime="00:04:48.90" resultid="6433" heatid="10945" lane="0" entrytime="00:04:43.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="100" swimtime="00:01:07.75" />
                    <SPLIT distance="150" swimtime="00:01:44.38" />
                    <SPLIT distance="200" swimtime="00:02:21.20" />
                    <SPLIT distance="250" swimtime="00:02:57.74" />
                    <SPLIT distance="300" swimtime="00:03:34.75" />
                    <SPLIT distance="350" swimtime="00:04:12.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WMT" nation="POL" region="14" clubid="5278" name="Warsaw Masters Team">
          <CONTACT city="Warszawa" email="wojciech.kaluzynski@gmail.com" name="Kałużyński Wojciech" phone="607 45 44444" state="MAZ" />
          <ATHLETES>
            <ATHLETE birthdate="1980-01-01" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="5534">
              <RESULTS>
                <RESULT eventid="1160" points="548" swimtime="00:00:25.54" resultid="8651" heatid="10710" lane="6" entrytime="00:00:25.00" />
                <RESULT eventid="1242" points="533" swimtime="00:00:29.65" resultid="8652" heatid="10751" lane="8" entrytime="00:00:29.80" />
                <RESULT eventid="1422" points="505" swimtime="00:00:28.15" resultid="8653" heatid="10826" lane="0" />
                <RESULT eventid="1452" points="487" swimtime="00:01:05.90" resultid="8654" heatid="10850" lane="6" entrytime="00:01:02.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="416" swimtime="00:02:29.90" resultid="8655" heatid="10899" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:13.67" />
                    <SPLIT distance="150" swimtime="00:01:52.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-16" firstname="Paweł" gender="M" lastname="Witkowski" nation="POL" athleteid="5421">
              <RESULTS>
                <RESULT eventid="1160" points="383" swimtime="00:00:28.79" resultid="8559" heatid="10699" lane="0" entrytime="00:00:31.50" />
                <RESULT eventid="1272" points="427" swimtime="00:02:48.62" resultid="8560" heatid="10762" lane="6" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:19.97" />
                    <SPLIT distance="150" swimtime="00:02:03.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="455" swimtime="00:01:14.25" resultid="8561" heatid="10817" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="519" swimtime="00:00:32.87" resultid="8562" heatid="10923" lane="0" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-04" firstname="Ewa" gender="F" lastname="Matlak" nation="POL" athleteid="5406">
              <RESULTS>
                <RESULT comment="G 8 - Ukończenie wyścigu nie w położeniu na plecach" eventid="1175" status="DSQ" swimtime="00:03:11.69" resultid="8547" heatid="10715" lane="6" entrytime="00:03:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:01:28.80" />
                    <SPLIT distance="150" swimtime="00:02:26.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="320" swimtime="00:01:16.08" resultid="8548" heatid="10770" lane="8" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="330" swimtime="00:00:35.33" resultid="8549" heatid="10822" lane="6" entrytime="00:00:37.80" />
                <RESULT eventid="1467" points="334" swimtime="00:02:42.82" resultid="8550" heatid="10854" lane="2" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:17.39" />
                    <SPLIT distance="150" swimtime="00:02:00.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="313" swimtime="00:05:48.17" resultid="8551" heatid="10934" lane="9" entrytime="00:05:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                    <SPLIT distance="100" swimtime="00:01:20.34" />
                    <SPLIT distance="150" swimtime="00:02:04.68" />
                    <SPLIT distance="200" swimtime="00:02:49.58" />
                    <SPLIT distance="250" swimtime="00:03:34.52" />
                    <SPLIT distance="300" swimtime="00:04:20.24" />
                    <SPLIT distance="350" swimtime="00:05:05.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-20" firstname="Katarzyna" gender="F" lastname="Dziedzic" nation="POL" athleteid="5546">
              <RESULTS>
                <RESULT eventid="1175" points="275" swimtime="00:03:13.93" resultid="8661" heatid="10716" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:01:29.43" />
                    <SPLIT distance="150" swimtime="00:02:25.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="277" swimtime="00:01:38.62" resultid="8662" heatid="10806" lane="7" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="266" swimtime="00:00:37.96" resultid="8663" heatid="10823" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1623" points="327" swimtime="00:00:42.78" resultid="8664" heatid="10909" lane="1" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-14" firstname="Sebastian" gender="M" lastname="Wojciechowski" nation="POL" athleteid="5309">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="8465" heatid="10693" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="8466" heatid="10777" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="8467" heatid="10860" lane="9" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="5347">
              <RESULTS>
                <RESULT eventid="1160" points="183" swimtime="00:00:36.82" resultid="8497" heatid="10693" lane="4" entrytime="00:00:37.03" />
                <RESULT eventid="1272" points="233" swimtime="00:03:26.37" resultid="8498" heatid="10759" lane="4" entrytime="00:03:26.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                    <SPLIT distance="100" swimtime="00:01:36.44" />
                    <SPLIT distance="150" swimtime="00:02:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="116" swimtime="00:03:48.30" resultid="8499" heatid="10792" lane="6" entrytime="00:03:58.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.61" />
                    <SPLIT distance="100" swimtime="00:01:48.90" />
                    <SPLIT distance="150" swimtime="00:02:49.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="222" swimtime="00:01:34.34" resultid="8500" heatid="10812" lane="3" entrytime="00:01:35.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="121" swimtime="00:01:40.56" resultid="8501" heatid="10886" lane="3" entrytime="00:01:36.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="262" swimtime="00:00:41.26" resultid="8502" heatid="10916" lane="7" entrytime="00:00:42.83" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="5412">
              <RESULTS>
                <RESULT eventid="1160" points="480" swimtime="00:00:26.70" resultid="8552" heatid="10709" lane="5" entrytime="00:00:25.90" />
                <RESULT eventid="1302" points="508" swimtime="00:00:58.77" resultid="8553" heatid="10787" lane="2" entrytime="00:00:57.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="504" swimtime="00:02:08.15" resultid="8554" heatid="10866" lane="8" entrytime="00:02:07.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="100" swimtime="00:01:01.89" />
                    <SPLIT distance="150" swimtime="00:01:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="470" swimtime="00:04:42.85" resultid="8555" heatid="10944" lane="1" entrytime="00:04:51.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:01:04.86" />
                    <SPLIT distance="150" swimtime="00:01:41.47" />
                    <SPLIT distance="200" swimtime="00:02:18.36" />
                    <SPLIT distance="250" swimtime="00:02:55.21" />
                    <SPLIT distance="300" swimtime="00:03:31.89" />
                    <SPLIT distance="350" swimtime="00:04:08.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisław" gender="M" lastname="Kozak" nation="POL" athleteid="5473">
              <RESULTS>
                <RESULT eventid="1160" points="272" swimtime="00:00:32.24" resultid="8602" heatid="10698" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1272" points="480" swimtime="00:02:42.21" resultid="8603" heatid="10764" lane="9" entrytime="00:02:42.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="500" swimtime="00:01:11.94" resultid="8604" heatid="10819" lane="2" entrytime="00:01:10.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="583" swimtime="00:00:31.61" resultid="8605" heatid="10926" lane="9" entrytime="00:00:31.77" />
                <RESULT eventid="1695" points="317" swimtime="00:05:22.53" resultid="9530" heatid="10943" lane="2" entrytime="00:05:03.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                    <SPLIT distance="150" swimtime="00:01:53.39" />
                    <SPLIT distance="200" swimtime="00:02:34.81" />
                    <SPLIT distance="250" swimtime="00:03:16.32" />
                    <SPLIT distance="300" swimtime="00:03:58.28" />
                    <SPLIT distance="350" swimtime="00:04:40.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-30" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="5386">
              <RESULTS>
                <RESULT eventid="1190" points="303" swimtime="00:02:49.56" resultid="8531" heatid="10725" lane="3" entrytime="00:02:49.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:01:17.43" />
                    <SPLIT distance="150" swimtime="00:02:11.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="375" swimtime="00:01:05.03" resultid="8532" heatid="10779" lane="3" entrytime="00:01:09.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="318" swimtime="00:01:15.96" resultid="8533" heatid="10843" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="339" swimtime="00:02:26.15" resultid="8534" heatid="10862" lane="1" entrytime="00:02:26.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:11.15" />
                    <SPLIT distance="150" swimtime="00:01:49.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="315" swimtime="00:02:44.39" resultid="8535" heatid="10902" lane="6" entrytime="00:02:48.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:01:19.14" />
                    <SPLIT distance="150" swimtime="00:02:01.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="5354">
              <RESULTS>
                <RESULT eventid="1160" points="436" swimtime="00:00:27.57" resultid="8503" heatid="10707" lane="9" entrytime="00:00:27.34" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  w  kat G  55-59  lat" eventid="1190" points="412" swimtime="00:02:33.14" resultid="8504" heatid="10728" lane="0" entrytime="00:02:36.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                    <SPLIT distance="150" swimtime="00:01:58.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="497" swimtime="00:00:59.19" resultid="8505" heatid="10785" lane="4" entrytime="00:00:59.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="396" swimtime="00:00:30.53" resultid="8506" heatid="10834" lane="0" entrytime="00:00:30.42" />
                <RESULT eventid="1482" points="443" swimtime="00:02:13.74" resultid="8507" heatid="10864" lane="4" entrytime="00:02:14.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:06.53" />
                    <SPLIT distance="150" swimtime="00:01:40.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="8508" heatid="10923" lane="8" entrytime="00:00:35.41" />
                <RESULT eventid="1695" points="430" swimtime="00:04:51.55" resultid="8509" heatid="10944" lane="8" entrytime="00:04:55.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                    <SPLIT distance="150" swimtime="00:01:49.50" />
                    <SPLIT distance="200" swimtime="00:02:26.78" />
                    <SPLIT distance="250" swimtime="00:03:03.72" />
                    <SPLIT distance="300" swimtime="00:03:40.14" />
                    <SPLIT distance="350" swimtime="00:04:16.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-12-04" firstname="Jacek" gender="M" lastname="Nowakowski" nation="POL" athleteid="5392">
              <RESULTS>
                <RESULT eventid="1128" points="259" swimtime="00:22:44.85" resultid="8536" heatid="10678" lane="8" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:20.70" />
                    <SPLIT distance="150" swimtime="00:02:05.52" />
                    <SPLIT distance="200" swimtime="00:02:50.96" />
                    <SPLIT distance="250" swimtime="00:03:36.98" />
                    <SPLIT distance="300" swimtime="00:04:22.51" />
                    <SPLIT distance="350" swimtime="00:05:08.78" />
                    <SPLIT distance="400" swimtime="00:05:54.60" />
                    <SPLIT distance="450" swimtime="00:06:40.59" />
                    <SPLIT distance="500" swimtime="00:07:26.75" />
                    <SPLIT distance="550" swimtime="00:08:12.61" />
                    <SPLIT distance="600" swimtime="00:08:58.66" />
                    <SPLIT distance="650" swimtime="00:09:44.44" />
                    <SPLIT distance="700" swimtime="00:10:30.72" />
                    <SPLIT distance="750" swimtime="00:11:17.05" />
                    <SPLIT distance="800" swimtime="00:12:03.31" />
                    <SPLIT distance="850" swimtime="00:12:48.95" />
                    <SPLIT distance="900" swimtime="00:13:35.20" />
                    <SPLIT distance="950" swimtime="00:14:21.16" />
                    <SPLIT distance="1000" swimtime="00:15:07.13" />
                    <SPLIT distance="1050" swimtime="00:15:53.33" />
                    <SPLIT distance="1100" swimtime="00:16:39.05" />
                    <SPLIT distance="1150" swimtime="00:17:24.88" />
                    <SPLIT distance="1200" swimtime="00:18:10.47" />
                    <SPLIT distance="1250" swimtime="00:18:56.31" />
                    <SPLIT distance="1300" swimtime="00:19:42.55" />
                    <SPLIT distance="1350" swimtime="00:20:27.89" />
                    <SPLIT distance="1400" swimtime="00:21:14.30" />
                    <SPLIT distance="1450" swimtime="00:22:00.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="258" swimtime="00:02:40.10" resultid="8537" heatid="10859" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:16.79" />
                    <SPLIT distance="150" swimtime="00:02:00.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="262" swimtime="00:05:43.54" resultid="8538" heatid="10940" lane="2" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:01.37" />
                    <SPLIT distance="200" swimtime="00:02:45.67" />
                    <SPLIT distance="250" swimtime="00:03:30.19" />
                    <SPLIT distance="300" swimtime="00:04:15.37" />
                    <SPLIT distance="350" swimtime="00:05:00.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-11-10" firstname="Anna" gender="F" lastname="Turczyn" nation="POL" athleteid="5329">
              <RESULTS>
                <RESULT eventid="1175" points="160" swimtime="00:03:51.89" resultid="8482" heatid="10713" lane="5" entrytime="00:03:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.33" />
                    <SPLIT distance="100" swimtime="00:01:59.72" />
                    <SPLIT distance="150" swimtime="00:02:57.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="238" swimtime="00:03:44.25" resultid="8483" heatid="10754" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.56" />
                    <SPLIT distance="100" swimtime="00:01:46.88" />
                    <SPLIT distance="150" swimtime="00:02:45.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="233" swimtime="00:01:44.51" resultid="8484" heatid="10805" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" status="DNS" swimtime="00:00:00.00" resultid="8485" heatid="10907" lane="6" entrytime="00:00:48.00" />
                <RESULT eventid="1674" points="189" swimtime="00:06:51.74" resultid="8486" heatid="10932" lane="2" entrytime="00:06:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.08" />
                    <SPLIT distance="100" swimtime="00:01:34.82" />
                    <SPLIT distance="150" swimtime="00:02:27.15" />
                    <SPLIT distance="200" swimtime="00:03:20.20" />
                    <SPLIT distance="250" swimtime="00:04:13.50" />
                    <SPLIT distance="300" swimtime="00:05:07.41" />
                    <SPLIT distance="350" swimtime="00:06:00.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-13" firstname="Agnieszka" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="5522">
              <RESULTS>
                <RESULT eventid="1287" points="277" swimtime="00:01:19.83" resultid="8641" heatid="10768" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="247" swimtime="00:02:59.84" resultid="8642" heatid="10853" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="100" swimtime="00:01:24.38" />
                    <SPLIT distance="150" swimtime="00:02:12.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="231" swimtime="00:06:25.13" resultid="8643" heatid="10932" lane="4" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                    <SPLIT distance="100" swimtime="00:01:32.60" />
                    <SPLIT distance="150" swimtime="00:02:22.19" />
                    <SPLIT distance="200" swimtime="00:03:12.93" />
                    <SPLIT distance="250" swimtime="00:04:01.66" />
                    <SPLIT distance="300" swimtime="00:04:50.43" />
                    <SPLIT distance="350" swimtime="00:05:38.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-20" firstname="Magdalena" gender="F" lastname="Mostowska" nation="POL" athleteid="5344">
              <RESULTS>
                <RESULT eventid="1113" points="233" swimtime="00:25:03.50" resultid="8495" heatid="10674" lane="1" entrytime="00:28:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.55" />
                    <SPLIT distance="100" swimtime="00:01:34.28" />
                    <SPLIT distance="150" swimtime="00:02:22.47" />
                    <SPLIT distance="200" swimtime="00:03:11.25" />
                    <SPLIT distance="250" swimtime="00:04:00.84" />
                    <SPLIT distance="300" swimtime="00:04:50.19" />
                    <SPLIT distance="350" swimtime="00:05:40.10" />
                    <SPLIT distance="400" swimtime="00:06:29.96" />
                    <SPLIT distance="450" swimtime="00:07:20.35" />
                    <SPLIT distance="500" swimtime="00:08:10.62" />
                    <SPLIT distance="550" swimtime="00:09:00.68" />
                    <SPLIT distance="600" swimtime="00:09:50.78" />
                    <SPLIT distance="650" swimtime="00:10:41.22" />
                    <SPLIT distance="700" swimtime="00:11:31.41" />
                    <SPLIT distance="750" swimtime="00:12:21.67" />
                    <SPLIT distance="800" swimtime="00:13:12.11" />
                    <SPLIT distance="850" swimtime="00:14:02.89" />
                    <SPLIT distance="900" swimtime="00:14:53.45" />
                    <SPLIT distance="950" swimtime="00:15:44.38" />
                    <SPLIT distance="1000" swimtime="00:16:35.32" />
                    <SPLIT distance="1050" swimtime="00:17:26.64" />
                    <SPLIT distance="1100" swimtime="00:18:17.88" />
                    <SPLIT distance="1150" swimtime="00:19:08.76" />
                    <SPLIT distance="1200" swimtime="00:19:59.58" />
                    <SPLIT distance="1250" swimtime="00:20:50.99" />
                    <SPLIT distance="1300" swimtime="00:21:41.93" />
                    <SPLIT distance="1350" swimtime="00:22:32.79" />
                    <SPLIT distance="1400" swimtime="00:23:23.78" />
                    <SPLIT distance="1450" swimtime="00:24:14.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="237" swimtime="00:06:21.77" resultid="8496" heatid="10932" lane="5" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                    <SPLIT distance="100" swimtime="00:01:31.03" />
                    <SPLIT distance="150" swimtime="00:02:18.73" />
                    <SPLIT distance="200" swimtime="00:03:06.88" />
                    <SPLIT distance="250" swimtime="00:03:55.69" />
                    <SPLIT distance="300" swimtime="00:04:44.69" />
                    <SPLIT distance="350" swimtime="00:05:34.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-10" firstname="Damian" gender="M" lastname="Rajzer" nation="POL" athleteid="5492">
              <RESULTS>
                <RESULT eventid="1160" points="356" swimtime="00:00:29.49" resultid="8617" heatid="10702" lane="9" entrytime="00:00:29.50" />
                <RESULT eventid="1302" points="318" swimtime="00:01:08.72" resultid="8618" heatid="10777" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNF" swimtime="00:00:00.00" resultid="8619" heatid="10833" lane="9" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-10" firstname="Katarzyna" gender="F" lastname="Czarnecka" nation="POL" athleteid="5483">
              <RESULTS>
                <RESULT eventid="1144" points="413" swimtime="00:00:31.84" resultid="8610" heatid="10686" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1257" points="294" swimtime="00:03:29.07" resultid="8611" heatid="10755" lane="0" entrytime="00:03:25.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.86" />
                    <SPLIT distance="100" swimtime="00:01:41.26" />
                    <SPLIT distance="150" swimtime="00:02:35.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="347" swimtime="00:01:31.52" resultid="8612" heatid="10807" lane="1" entrytime="00:01:30.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="399" swimtime="00:00:40.02" resultid="8613" heatid="10910" lane="6" entrytime="00:00:39.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-13" firstname="Marcin" gender="M" lastname="Giejsztowt" nation="POL" athleteid="5438">
              <RESULTS>
                <RESULT eventid="1128" points="387" swimtime="00:19:55.11" resultid="8573" heatid="10679" lane="0" entrytime="00:20:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:49.50" />
                    <SPLIT distance="200" swimtime="00:02:29.63" />
                    <SPLIT distance="250" swimtime="00:03:10.06" />
                    <SPLIT distance="300" swimtime="00:03:50.31" />
                    <SPLIT distance="350" swimtime="00:04:30.49" />
                    <SPLIT distance="400" swimtime="00:05:10.85" />
                    <SPLIT distance="450" swimtime="00:05:50.93" />
                    <SPLIT distance="500" swimtime="00:06:31.91" />
                    <SPLIT distance="550" swimtime="00:07:12.31" />
                    <SPLIT distance="600" swimtime="00:07:53.14" />
                    <SPLIT distance="650" swimtime="00:08:33.57" />
                    <SPLIT distance="700" swimtime="00:09:15.14" />
                    <SPLIT distance="750" swimtime="00:09:55.48" />
                    <SPLIT distance="800" swimtime="00:10:35.84" />
                    <SPLIT distance="850" swimtime="00:11:15.86" />
                    <SPLIT distance="900" swimtime="00:11:56.39" />
                    <SPLIT distance="950" swimtime="00:12:36.58" />
                    <SPLIT distance="1000" swimtime="00:13:17.51" />
                    <SPLIT distance="1050" swimtime="00:13:57.29" />
                    <SPLIT distance="1100" swimtime="00:14:38.22" />
                    <SPLIT distance="1150" swimtime="00:15:18.11" />
                    <SPLIT distance="1200" swimtime="00:15:59.32" />
                    <SPLIT distance="1250" swimtime="00:16:38.95" />
                    <SPLIT distance="1300" swimtime="00:17:19.76" />
                    <SPLIT distance="1350" swimtime="00:17:59.75" />
                    <SPLIT distance="1400" swimtime="00:18:40.52" />
                    <SPLIT distance="1450" swimtime="00:19:19.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="413" swimtime="00:01:02.95" resultid="8574" heatid="10782" lane="0" entrytime="00:01:04.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="411" swimtime="00:02:17.17" resultid="8575" heatid="10862" lane="3" entrytime="00:02:22.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:05.80" />
                    <SPLIT distance="150" swimtime="00:01:41.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="402" swimtime="00:04:58.03" resultid="8576" heatid="10943" lane="4" entrytime="00:05:02.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:49.32" />
                    <SPLIT distance="200" swimtime="00:02:27.62" />
                    <SPLIT distance="250" swimtime="00:03:05.36" />
                    <SPLIT distance="300" swimtime="00:03:43.80" />
                    <SPLIT distance="350" swimtime="00:04:21.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-04-14" firstname="Wiesław" gender="M" lastname="Załuski" nation="POL" athleteid="5300">
              <RESULTS>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="8458" heatid="10723" lane="2" entrytime="00:03:02.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn w  kat I  65-69  lat" eventid="1242" points="277" swimtime="00:00:36.86" resultid="8459" heatid="10746" lane="6" entrytime="00:00:37.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Mężczyzn  w  kat I  65-69  lat" eventid="1452" points="240" swimtime="00:01:23.33" resultid="8460" heatid="10847" lane="0" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1608" points="199" swimtime="00:03:11.66" resultid="8461" heatid="10902" lane="9" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.54" />
                    <SPLIT distance="100" swimtime="00:01:32.92" />
                    <SPLIT distance="150" swimtime="00:02:22.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="5313">
              <RESULTS>
                <RESULT eventid="1160" points="487" swimtime="00:00:26.57" resultid="8468" heatid="10706" lane="6" entrytime="00:00:27.50" />
                <RESULT eventid="1302" points="577" swimtime="00:00:56.33" resultid="8469" heatid="10785" lane="0" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="594" swimtime="00:00:26.68" resultid="8470" heatid="10838" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="1546" status="DNS" swimtime="00:00:00.00" resultid="8471" heatid="10880" lane="3" entrytime="00:05:30.00" />
                <RESULT eventid="1578" points="498" swimtime="00:01:02.85" resultid="8472" heatid="10892" lane="7" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 14 - Praca nóg  w płaszczyźnie pionowej w dół /z wyjątkiem jednego ruchu po starcie i nawrocie/" eventid="1638" status="DSQ" swimtime="00:00:34.15" resultid="8473" heatid="10923" lane="7" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-05" firstname="Bartłomiej" gender="M" lastname="Pawłowski" nation="POL" athleteid="5462">
              <RESULTS>
                <RESULT eventid="1160" points="345" swimtime="00:00:29.81" resultid="8593" heatid="10702" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1302" points="332" swimtime="00:01:07.69" resultid="8594" heatid="10781" lane="9" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="295" swimtime="00:01:25.74" resultid="8595" heatid="10815" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="391" swimtime="00:00:36.13" resultid="8596" heatid="10921" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-05-15" firstname="Jerzy" gender="M" lastname="Leszczyński" nation="POL" athleteid="5467">
              <RESULTS>
                <RESULT eventid="1160" points="335" swimtime="00:00:30.08" resultid="8597" heatid="10701" lane="6" entrytime="00:00:29.80" />
                <RESULT eventid="1190" points="268" swimtime="00:02:56.68" resultid="8598" heatid="10724" lane="5" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:24.87" />
                    <SPLIT distance="150" swimtime="00:02:15.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="273" swimtime="00:03:15.68" resultid="8599" heatid="10761" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                    <SPLIT distance="100" swimtime="00:01:31.61" />
                    <SPLIT distance="150" swimtime="00:02:23.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="301" swimtime="00:01:09.97" resultid="8600" heatid="10780" lane="0" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="277" swimtime="00:01:27.63" resultid="8601" heatid="10815" lane="8" entrytime="00:01:25.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-09-27" firstname="Wojciech" gender="M" lastname="Kossowski" nation="POL" athleteid="5417">
              <RESULTS>
                <RESULT eventid="1190" points="162" swimtime="00:03:28.89" resultid="8556" heatid="10721" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                    <SPLIT distance="100" swimtime="00:01:44.28" />
                    <SPLIT distance="150" swimtime="00:02:41.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="194" swimtime="00:03:39.28" resultid="8557" heatid="10760" lane="0" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.57" />
                    <SPLIT distance="100" swimtime="00:01:41.44" />
                    <SPLIT distance="150" swimtime="00:02:39.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="223" swimtime="00:01:34.19" resultid="8558" heatid="10813" lane="7" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-11-24" firstname="Krzysztof" gender="M" lastname="Gogol" nation="POL" athleteid="5296">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="8455" heatid="10694" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="8456" heatid="10776" lane="8" entrytime="00:01:20.00" />
                <RESULT eventid="1482" status="DNS" swimtime="00:00:00.00" resultid="8457" heatid="10856" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-10-11" firstname="Grzegorz" gender="M" lastname="Matyszewski" nation="POL" athleteid="5320">
              <RESULTS>
                <RESULT eventid="1160" points="265" swimtime="00:00:32.55" resultid="8474" heatid="10695" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1190" points="193" swimtime="00:03:17.02" resultid="8475" heatid="10721" lane="5" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                    <SPLIT distance="100" swimtime="00:01:35.77" />
                    <SPLIT distance="150" swimtime="00:02:30.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="255" swimtime="00:03:20.17" resultid="8476" heatid="10759" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                    <SPLIT distance="100" swimtime="00:01:33.59" />
                    <SPLIT distance="150" swimtime="00:02:26.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="220" swimtime="00:01:17.68" resultid="8477" heatid="10776" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="273" swimtime="00:01:28.00" resultid="8478" heatid="10814" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="168" swimtime="00:03:04.63" resultid="8479" heatid="10858" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:27.98" />
                    <SPLIT distance="150" swimtime="00:02:17.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="311" swimtime="00:00:38.99" resultid="8480" heatid="10919" lane="7" entrytime="00:00:39.15" />
                <RESULT eventid="1695" points="144" swimtime="00:06:59.55" resultid="8481" heatid="10937" lane="1" entrytime="00:06:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                    <SPLIT distance="100" swimtime="00:01:31.74" />
                    <SPLIT distance="150" swimtime="00:02:24.75" />
                    <SPLIT distance="200" swimtime="00:03:18.30" />
                    <SPLIT distance="250" swimtime="00:04:13.09" />
                    <SPLIT distance="300" swimtime="00:05:08.35" />
                    <SPLIT distance="350" swimtime="00:06:05.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-13" firstname="Rafał" gender="M" lastname="Tichy" nation="POL" athleteid="5488">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="8614" heatid="10694" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="8615" heatid="10775" lane="8" entrytime="00:01:25.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="8616" heatid="10827" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-11-11" firstname="Bolesław" gender="M" lastname="Szuter" nation="POL" athleteid="5396">
              <RESULTS>
                <RESULT eventid="1160" points="500" swimtime="00:00:26.34" resultid="8539" heatid="10709" lane="4" entrytime="00:00:25.79" />
                <RESULT eventid="1302" points="575" swimtime="00:00:56.39" resultid="8540" heatid="10788" lane="9" entrytime="00:00:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="524" swimtime="00:02:06.51" resultid="8541" heatid="10866" lane="2" entrytime="00:02:04.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="100" swimtime="00:01:02.13" />
                    <SPLIT distance="150" swimtime="00:01:34.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Mężczyzn w  kat E  45-49  lat" eventid="1422" points="519" swimtime="00:00:27.90" resultid="9051" heatid="10836" lane="5" entrytime="00:00:28.23" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="5400">
              <RESULTS>
                <RESULT eventid="1190" points="43" swimtime="00:05:23.19" resultid="8542" heatid="10719" lane="2" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.41" />
                    <SPLIT distance="100" swimtime="00:02:41.03" />
                    <SPLIT distance="150" swimtime="00:04:08.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="8543" heatid="10740" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="8544" heatid="10809" lane="5" entrytime="00:02:45.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="8545" heatid="10826" lane="7" entrytime="00:01:25.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="8546" heatid="10913" lane="8" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-06-10" firstname="Łukasz" gender="M" lastname="Rybiński" nation="POL" athleteid="5335">
              <RESULTS>
                <RESULT eventid="1160" points="320" swimtime="00:00:30.57" resultid="8487" heatid="10700" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="8488" heatid="10722" lane="6" entrytime="00:03:10.00" />
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="8489" heatid="10745" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1302" points="307" swimtime="00:01:09.52" resultid="8490" heatid="10779" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="268" swimtime="00:01:28.52" resultid="8491" heatid="10814" lane="8" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="8492" heatid="10828" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1638" points="305" swimtime="00:00:39.24" resultid="8493" heatid="10919" lane="8" entrytime="00:00:39.50" />
                <RESULT eventid="1695" points="215" swimtime="00:06:06.99" resultid="8494" heatid="10939" lane="6" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                    <SPLIT distance="100" swimtime="00:01:20.45" />
                    <SPLIT distance="150" swimtime="00:02:05.69" />
                    <SPLIT distance="200" swimtime="00:02:52.85" />
                    <SPLIT distance="250" swimtime="00:03:40.60" />
                    <SPLIT distance="300" swimtime="00:04:29.75" />
                    <SPLIT distance="350" swimtime="00:05:19.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka - Skorykow" nation="POL" athleteid="5518">
              <RESULTS>
                <RESULT eventid="1144" points="394" swimtime="00:00:32.36" resultid="9487" heatid="10686" lane="0" entrytime="00:00:33.50" />
                <RESULT eventid="1376" points="330" swimtime="00:01:33.06" resultid="9488" heatid="10806" lane="0" entrytime="00:01:39.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="370" swimtime="00:00:41.03" resultid="9489" heatid="10909" lane="0" entrytime="00:00:43.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michał" gender="M" lastname="Nowak" nation="POL" athleteid="5509">
              <RESULTS>
                <RESULT eventid="1190" points="224" swimtime="00:03:07.44" resultid="8631" heatid="10722" lane="5" entrytime="00:03:09.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                    <SPLIT distance="100" swimtime="00:01:32.47" />
                    <SPLIT distance="150" swimtime="00:02:22.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="269" swimtime="00:03:16.72" resultid="8632" heatid="10760" lane="4" entrytime="00:03:15.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                    <SPLIT distance="100" swimtime="00:01:32.83" />
                    <SPLIT distance="150" swimtime="00:02:24.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="292" swimtime="00:01:26.09" resultid="8633" heatid="10815" lane="0" entrytime="00:01:26.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="189" swimtime="00:07:04.22" resultid="8634" heatid="10877" lane="6" entrytime="00:07:09.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.78" />
                    <SPLIT distance="100" swimtime="00:01:52.50" />
                    <SPLIT distance="150" swimtime="00:02:48.43" />
                    <SPLIT distance="200" swimtime="00:03:44.28" />
                    <SPLIT distance="250" swimtime="00:04:38.61" />
                    <SPLIT distance="300" swimtime="00:05:32.96" />
                    <SPLIT distance="350" swimtime="00:06:19.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="354" swimtime="00:00:37.32" resultid="8635" heatid="10920" lane="1" entrytime="00:00:38.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-07-10" firstname="Daniel" gender="M" lastname="Julian" nation="POL" athleteid="5279">
              <RESULTS>
                <RESULT eventid="1098" points="372" swimtime="00:10:28.46" resultid="8440" heatid="10671" lane="3" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:51.02" />
                    <SPLIT distance="200" swimtime="00:02:31.49" />
                    <SPLIT distance="250" swimtime="00:03:11.55" />
                    <SPLIT distance="300" swimtime="00:03:52.01" />
                    <SPLIT distance="350" swimtime="00:04:32.32" />
                    <SPLIT distance="400" swimtime="00:05:12.45" />
                    <SPLIT distance="450" swimtime="00:05:52.69" />
                    <SPLIT distance="500" swimtime="00:06:33.14" />
                    <SPLIT distance="550" swimtime="00:07:13.66" />
                    <SPLIT distance="600" swimtime="00:07:53.57" />
                    <SPLIT distance="650" swimtime="00:08:33.17" />
                    <SPLIT distance="700" swimtime="00:09:12.65" />
                    <SPLIT distance="750" swimtime="00:09:51.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="481" swimtime="00:00:26.68" resultid="8441" heatid="10706" lane="8" entrytime="00:00:27.50" />
                <RESULT eventid="1242" points="443" swimtime="00:00:31.52" resultid="8442" heatid="10750" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1302" points="504" swimtime="00:00:58.94" resultid="8443" heatid="10786" lane="9" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="450" swimtime="00:01:07.62" resultid="8444" heatid="10849" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="434" swimtime="00:02:14.72" resultid="8445" heatid="10864" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:06.24" />
                    <SPLIT distance="150" swimtime="00:01:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="388" swimtime="00:02:33.40" resultid="8446" heatid="10903" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:15.30" />
                    <SPLIT distance="150" swimtime="00:01:55.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="421" swimtime="00:04:53.57" resultid="8447" heatid="10944" lane="9" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:08.60" />
                    <SPLIT distance="150" swimtime="00:01:45.80" />
                    <SPLIT distance="200" swimtime="00:02:23.47" />
                    <SPLIT distance="250" swimtime="00:03:01.45" />
                    <SPLIT distance="300" swimtime="00:03:39.08" />
                    <SPLIT distance="350" swimtime="00:04:16.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="5433">
              <RESULTS>
                <RESULT eventid="1059" points="108" swimtime="00:16:55.30" resultid="8569" heatid="10666" lane="7" entrytime="00:17:06.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.70" />
                    <SPLIT distance="100" swimtime="00:02:01.53" />
                    <SPLIT distance="150" swimtime="00:03:06.14" />
                    <SPLIT distance="200" swimtime="00:04:10.51" />
                    <SPLIT distance="250" swimtime="00:05:15.40" />
                    <SPLIT distance="300" swimtime="00:06:19.37" />
                    <SPLIT distance="350" swimtime="00:07:22.62" />
                    <SPLIT distance="400" swimtime="00:08:27.00" />
                    <SPLIT distance="450" swimtime="00:09:31.09" />
                    <SPLIT distance="500" swimtime="00:10:35.58" />
                    <SPLIT distance="550" swimtime="00:11:39.46" />
                    <SPLIT distance="600" swimtime="00:12:43.41" />
                    <SPLIT distance="650" swimtime="00:13:47.58" />
                    <SPLIT distance="700" swimtime="00:14:51.30" />
                    <SPLIT distance="750" swimtime="00:15:54.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="95" swimtime="00:00:51.88" resultid="8570" heatid="10681" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="1467" points="92" swimtime="00:04:09.56" resultid="8571" heatid="10851" lane="3" entrytime="00:04:10.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.00" />
                    <SPLIT distance="100" swimtime="00:01:59.39" />
                    <SPLIT distance="150" swimtime="00:03:06.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="98" swimtime="00:08:32.32" resultid="8572" heatid="10931" lane="1" entrytime="00:08:30.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.16" />
                    <SPLIT distance="100" swimtime="00:02:02.42" />
                    <SPLIT distance="150" swimtime="00:03:10.25" />
                    <SPLIT distance="200" swimtime="00:04:15.64" />
                    <SPLIT distance="250" swimtime="00:05:22.14" />
                    <SPLIT distance="300" swimtime="00:06:26.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-16" firstname="Tadeusz" gender="M" lastname="Vorbrodt" nation="POL" athleteid="5505">
              <RESULTS>
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="8628" heatid="10740" lane="2" />
                <RESULT eventid="1452" points="79" swimtime="00:02:00.56" resultid="8629" heatid="10844" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="122" swimtime="00:07:23.48" resultid="8630" heatid="10935" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:39.17" />
                    <SPLIT distance="150" swimtime="00:02:35.34" />
                    <SPLIT distance="200" swimtime="00:03:33.70" />
                    <SPLIT distance="250" swimtime="00:04:31.12" />
                    <SPLIT distance="300" swimtime="00:05:29.74" />
                    <SPLIT distance="350" swimtime="00:06:28.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-31" firstname="Katharina" gender="F" lastname="Szymańska" nation="POL" athleteid="5452">
              <RESULTS>
                <RESULT eventid="1593" points="124" swimtime="00:04:08.52" resultid="8585" heatid="10893" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.00" />
                    <SPLIT distance="100" swimtime="00:02:06.69" />
                    <SPLIT distance="150" swimtime="00:03:09.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1674" points="158" swimtime="00:07:16.73" resultid="8586" heatid="10930" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.92" />
                    <SPLIT distance="100" swimtime="00:01:46.31" />
                    <SPLIT distance="150" swimtime="00:02:42.36" />
                    <SPLIT distance="200" swimtime="00:03:38.60" />
                    <SPLIT distance="250" swimtime="00:04:34.27" />
                    <SPLIT distance="300" swimtime="00:05:30.74" />
                    <SPLIT distance="350" swimtime="00:06:27.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-21" firstname="Marianna" gender="F" lastname="Gajdus" nation="POL" athleteid="5540">
              <RESULTS>
                <RESULT eventid="1175" points="340" swimtime="00:03:00.63" resultid="9498" heatid="10716" lane="6" entrytime="00:03:01.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:26.74" />
                    <SPLIT distance="150" swimtime="00:02:19.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1317" points="246" swimtime="00:03:14.24" resultid="9499" heatid="10790" lane="6" entrytime="00:03:15.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:01:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="290" swimtime="00:01:37.17" resultid="9500" heatid="10806" lane="6" entrytime="00:01:35.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="303" swimtime="00:00:36.37" resultid="9501" heatid="10822" lane="4" entrytime="00:00:36.53" />
                <RESULT eventid="1562" points="296" swimtime="00:01:23.21" resultid="9502" heatid="10884" lane="8" entrytime="00:01:22.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="5371">
              <RESULTS>
                <RESULT eventid="1160" points="388" swimtime="00:00:28.65" resultid="8518" heatid="10700" lane="4" entrytime="00:00:30.01" />
                <RESULT eventid="1190" points="376" swimtime="00:02:37.81" resultid="8519" heatid="10727" lane="6" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:14.60" />
                    <SPLIT distance="150" swimtime="00:02:03.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="367" swimtime="00:00:33.57" resultid="8520" heatid="10749" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1302" points="444" swimtime="00:01:01.45" resultid="8521" heatid="10784" lane="1" entrytime="00:01:01.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="390" swimtime="00:01:10.96" resultid="8522" heatid="10849" lane="7" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="397" swimtime="00:02:18.67" resultid="8523" heatid="10863" lane="9" entrytime="00:02:20.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:08.56" />
                    <SPLIT distance="150" swimtime="00:01:43.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="348" swimtime="00:02:39.08" resultid="8524" heatid="10903" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:01:57.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-10-06" firstname="Mateusz" gender="M" lastname="Bednarz" nation="POL" athleteid="5455">
              <RESULTS>
                <RESULT eventid="1098" points="355" swimtime="00:10:37.97" resultid="8587" heatid="10672" lane="8" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="150" swimtime="00:01:50.74" />
                    <SPLIT distance="200" swimtime="00:02:29.93" />
                    <SPLIT distance="250" swimtime="00:03:10.21" />
                    <SPLIT distance="300" swimtime="00:03:49.79" />
                    <SPLIT distance="350" swimtime="00:04:30.76" />
                    <SPLIT distance="400" swimtime="00:05:10.86" />
                    <SPLIT distance="450" swimtime="00:05:51.77" />
                    <SPLIT distance="500" swimtime="00:06:32.51" />
                    <SPLIT distance="550" swimtime="00:07:13.83" />
                    <SPLIT distance="600" swimtime="00:07:54.47" />
                    <SPLIT distance="650" swimtime="00:08:35.60" />
                    <SPLIT distance="700" swimtime="00:09:17.70" />
                    <SPLIT distance="750" swimtime="00:09:59.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="338" swimtime="00:02:43.64" resultid="8588" heatid="10726" lane="7" entrytime="00:02:44.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                    <SPLIT distance="100" swimtime="00:01:19.50" />
                    <SPLIT distance="150" swimtime="00:02:07.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="8589" heatid="10746" lane="1" entrytime="00:00:37.27" />
                <RESULT eventid="1302" points="417" swimtime="00:01:02.77" resultid="8590" heatid="10782" lane="7" entrytime="00:01:03.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="406" swimtime="00:02:17.71" resultid="8591" heatid="10862" lane="4" entrytime="00:02:20.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:06.40" />
                    <SPLIT distance="150" swimtime="00:01:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="394" swimtime="00:05:00.09" resultid="8592" heatid="10942" lane="5" entrytime="00:05:08.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:11.64" />
                    <SPLIT distance="150" swimtime="00:01:49.81" />
                    <SPLIT distance="200" swimtime="00:02:28.93" />
                    <SPLIT distance="250" swimtime="00:03:07.73" />
                    <SPLIT distance="300" swimtime="00:03:46.08" />
                    <SPLIT distance="350" swimtime="00:04:24.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="5362">
              <RESULTS>
                <RESULT eventid="1098" points="152" swimtime="00:14:05.59" resultid="8510" heatid="10669" lane="4" entrytime="00:14:03.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.18" />
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                    <SPLIT distance="150" swimtime="00:02:32.86" />
                    <SPLIT distance="200" swimtime="00:03:26.11" />
                    <SPLIT distance="250" swimtime="00:04:19.62" />
                    <SPLIT distance="300" swimtime="00:05:13.41" />
                    <SPLIT distance="350" swimtime="00:06:06.23" />
                    <SPLIT distance="400" swimtime="00:06:59.58" />
                    <SPLIT distance="450" swimtime="00:07:53.41" />
                    <SPLIT distance="500" swimtime="00:08:46.55" />
                    <SPLIT distance="550" swimtime="00:09:40.29" />
                    <SPLIT distance="600" swimtime="00:10:34.88" />
                    <SPLIT distance="650" swimtime="00:11:29.29" />
                    <SPLIT distance="700" swimtime="00:12:22.91" />
                    <SPLIT distance="750" swimtime="00:13:15.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="148" swimtime="00:00:39.52" resultid="8511" heatid="10693" lane="0" entrytime="00:00:39.10" />
                <RESULT eventid="1242" points="83" swimtime="00:00:55.01" resultid="8512" heatid="10742" lane="0" entrytime="00:00:54.96" />
                <RESULT eventid="1302" points="165" swimtime="00:01:25.50" resultid="8513" heatid="10774" lane="3" entrytime="00:01:28.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="108" swimtime="00:00:46.99" resultid="8514" heatid="10827" lane="0" entrytime="00:00:46.76" />
                <RESULT eventid="1482" points="165" swimtime="00:03:05.81" resultid="8515" heatid="10858" lane="1" entrytime="00:03:09.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="100" swimtime="00:01:30.23" />
                    <SPLIT distance="150" swimtime="00:02:19.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="89" swimtime="00:01:51.31" resultid="8516" heatid="10885" lane="4" entrytime="00:01:58.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="168" swimtime="00:06:38.19" resultid="8517" heatid="10937" lane="2" entrytime="00:06:47.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                    <SPLIT distance="100" swimtime="00:01:34.61" />
                    <SPLIT distance="150" swimtime="00:02:25.70" />
                    <SPLIT distance="200" swimtime="00:03:17.66" />
                    <SPLIT distance="250" swimtime="00:04:08.91" />
                    <SPLIT distance="300" swimtime="00:04:59.91" />
                    <SPLIT distance="350" swimtime="00:05:51.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-06-07" firstname="Olga" gender="F" lastname="Krysiak" nation="POL" athleteid="5515">
              <RESULTS>
                <RESULT eventid="1144" points="530" swimtime="00:00:29.31" resultid="8636" heatid="10688" lane="1" entrytime="00:00:29.20" />
                <RESULT eventid="1287" points="507" swimtime="00:01:05.26" resultid="8637" heatid="10771" lane="7" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-22" firstname="Timea" gender="F" lastname="Balajcza" nation="POL" athleteid="5496">
              <RESULTS>
                <RESULT eventid="1144" points="265" swimtime="00:00:36.92" resultid="8620" heatid="10684" lane="6" entrytime="00:00:35.94" />
                <RESULT eventid="1175" points="246" swimtime="00:03:21.15" resultid="8621" heatid="10714" lane="3" entrytime="00:03:30.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:41.86" />
                    <SPLIT distance="150" swimtime="00:02:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="292" swimtime="00:03:29.54" resultid="8622" heatid="10755" lane="7" entrytime="00:03:24.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.26" />
                    <SPLIT distance="100" swimtime="00:01:41.82" />
                    <SPLIT distance="150" swimtime="00:02:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="219" swimtime="00:01:26.29" resultid="8623" heatid="10768" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="305" swimtime="00:01:35.51" resultid="8624" heatid="10807" lane="0" entrytime="00:01:33.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="229" swimtime="00:03:04.56" resultid="8625" heatid="10853" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                    <SPLIT distance="100" swimtime="00:01:28.34" />
                    <SPLIT distance="150" swimtime="00:02:16.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="317" swimtime="00:00:43.23" resultid="8627" heatid="10909" lane="7" entrytime="00:00:42.67" />
                <RESULT eventid="1674" points="218" swimtime="00:06:32.59" resultid="9373" heatid="10932" lane="3" entrytime="00:06:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:01:32.80" />
                    <SPLIT distance="200" swimtime="00:03:12.74" />
                    <SPLIT distance="250" swimtime="00:04:02.59" />
                    <SPLIT distance="300" swimtime="00:04:52.64" />
                    <SPLIT distance="350" swimtime="00:05:42.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="5526">
              <RESULTS>
                <RESULT eventid="1098" points="383" swimtime="00:10:22.14" resultid="8644" heatid="10673" lane="8" entrytime="00:10:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:13.90" />
                    <SPLIT distance="150" swimtime="00:01:53.16" />
                    <SPLIT distance="200" swimtime="00:02:31.95" />
                    <SPLIT distance="250" swimtime="00:03:10.95" />
                    <SPLIT distance="300" swimtime="00:03:50.23" />
                    <SPLIT distance="350" swimtime="00:04:29.70" />
                    <SPLIT distance="400" swimtime="00:05:08.98" />
                    <SPLIT distance="450" swimtime="00:05:48.18" />
                    <SPLIT distance="500" swimtime="00:06:27.29" />
                    <SPLIT distance="550" swimtime="00:07:07.33" />
                    <SPLIT distance="600" swimtime="00:07:46.65" />
                    <SPLIT distance="650" swimtime="00:08:26.00" />
                    <SPLIT distance="700" swimtime="00:09:05.28" />
                    <SPLIT distance="750" swimtime="00:09:44.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="439" swimtime="00:00:27.51" resultid="8645" heatid="10706" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="1242" points="413" swimtime="00:00:32.28" resultid="8646" heatid="10750" lane="9" entrytime="00:00:31.05" />
                <RESULT eventid="1332" status="DNS" swimtime="00:00:00.00" resultid="8647" heatid="10796" lane="0" entrytime="00:02:32.00" />
                <RESULT eventid="1422" points="453" swimtime="00:00:29.19" resultid="8648" heatid="10836" lane="1" entrytime="00:00:28.50" />
                <RESULT eventid="1482" points="386" swimtime="00:02:20.05" resultid="8649" heatid="10864" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:08.42" />
                    <SPLIT distance="150" swimtime="00:01:45.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="8650" heatid="10891" lane="2" entrytime="00:01:04.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-28" firstname="Paweł" gender="M" lastname="Rogosz" nation="POL" athleteid="5288">
              <RESULTS>
                <RESULT eventid="1160" points="363" swimtime="00:00:29.31" resultid="8448" heatid="10701" lane="3" entrytime="00:00:29.89" />
                <RESULT eventid="1190" points="384" swimtime="00:02:36.77" resultid="8449" heatid="10727" lane="7" entrytime="00:02:38.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:16.96" />
                    <SPLIT distance="150" swimtime="00:02:00.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="395" swimtime="00:02:53.00" resultid="8450" heatid="10762" lane="1" entrytime="00:02:59.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:02:07.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1332" points="286" swimtime="00:02:49.13" resultid="8451" heatid="10795" lane="8" entrytime="00:02:46.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:18.55" />
                    <SPLIT distance="150" swimtime="00:02:05.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1546" points="376" swimtime="00:05:37.56" resultid="8452" heatid="10880" lane="8" entrytime="00:05:46.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:20.77" />
                    <SPLIT distance="150" swimtime="00:02:05.48" />
                    <SPLIT distance="200" swimtime="00:02:51.53" />
                    <SPLIT distance="250" swimtime="00:03:37.29" />
                    <SPLIT distance="300" swimtime="00:04:23.34" />
                    <SPLIT distance="350" swimtime="00:05:00.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="8453" heatid="10889" lane="0" entrytime="00:01:14.25" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="8454" heatid="10923" lane="9" entrytime="00:00:35.78" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="Borodziuk" nation="POL" athleteid="5443">
              <RESULTS>
                <RESULT eventid="1098" points="87" swimtime="00:17:00.13" resultid="8577" heatid="10669" lane="5" entrytime="00:16:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.05" />
                    <SPLIT distance="100" swimtime="00:01:50.12" />
                    <SPLIT distance="150" swimtime="00:02:51.58" />
                    <SPLIT distance="200" swimtime="00:03:58.89" />
                    <SPLIT distance="250" swimtime="00:05:04.59" />
                    <SPLIT distance="300" swimtime="00:06:09.69" />
                    <SPLIT distance="350" swimtime="00:07:16.10" />
                    <SPLIT distance="400" swimtime="00:08:24.20" />
                    <SPLIT distance="450" swimtime="00:09:27.64" />
                    <SPLIT distance="500" swimtime="00:10:35.77" />
                    <SPLIT distance="550" swimtime="00:11:40.40" />
                    <SPLIT distance="600" swimtime="00:12:48.59" />
                    <SPLIT distance="650" swimtime="00:13:53.19" />
                    <SPLIT distance="700" swimtime="00:14:59.90" />
                    <SPLIT distance="750" swimtime="00:16:05.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="173" swimtime="00:00:37.50" resultid="8578" heatid="10693" lane="3" entrytime="00:00:37.50" />
                <RESULT eventid="1242" points="113" swimtime="00:00:49.68" resultid="8579" heatid="10742" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1302" points="151" swimtime="00:01:28.04" resultid="8580" heatid="10774" lane="4" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="85" swimtime="00:01:57.91" resultid="8581" heatid="10845" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="85" swimtime="00:03:51.42" resultid="8582" heatid="10857" lane="5" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.87" />
                    <SPLIT distance="100" swimtime="00:01:45.99" />
                    <SPLIT distance="150" swimtime="00:02:51.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="8583" heatid="10900" lane="0" entrytime="00:04:10.00" />
                <RESULT eventid="1695" points="97" swimtime="00:07:57.85" resultid="8584" heatid="10936" lane="4" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.68" />
                    <SPLIT distance="100" swimtime="00:01:50.33" />
                    <SPLIT distance="150" swimtime="00:02:53.63" />
                    <SPLIT distance="200" swimtime="00:03:56.94" />
                    <SPLIT distance="250" swimtime="00:05:00.79" />
                    <SPLIT distance="300" swimtime="00:06:02.94" />
                    <SPLIT distance="350" swimtime="00:07:04.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-13" firstname="Michał" gender="M" lastname="Jabłoński" nation="POL" athleteid="5379">
              <RESULTS>
                <RESULT eventid="1160" points="353" swimtime="00:00:29.56" resultid="8525" heatid="10701" lane="5" entrytime="00:00:29.76" />
                <RESULT eventid="1302" points="367" swimtime="00:01:05.50" resultid="8526" heatid="10780" lane="6" entrytime="00:01:06.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="364" swimtime="00:00:31.40" resultid="8527" heatid="10832" lane="0" entrytime="00:00:32.40" />
                <RESULT eventid="1482" points="327" swimtime="00:02:28.00" resultid="8528" heatid="10861" lane="4" entrytime="00:02:28.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:11.18" />
                    <SPLIT distance="150" swimtime="00:01:49.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="320" swimtime="00:01:12.83" resultid="8529" heatid="10888" lane="2" entrytime="00:01:17.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="325" swimtime="00:05:19.84" resultid="8530" heatid="10941" lane="6" entrytime="00:05:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:14.83" />
                    <SPLIT distance="150" swimtime="00:01:55.58" />
                    <SPLIT distance="200" swimtime="00:02:36.93" />
                    <SPLIT distance="250" swimtime="00:03:18.03" />
                    <SPLIT distance="300" swimtime="00:03:59.09" />
                    <SPLIT distance="350" swimtime="00:04:40.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-14" firstname="Bartosz" gender="M" lastname="Ostrowski" nation="POL" athleteid="5426">
              <RESULTS>
                <RESULT eventid="1190" points="273" swimtime="00:02:55.71" resultid="8563" heatid="10723" lane="0" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                    <SPLIT distance="100" swimtime="00:01:27.10" />
                    <SPLIT distance="150" swimtime="00:02:15.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="274" swimtime="00:00:36.97" resultid="8564" heatid="10745" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1302" points="346" swimtime="00:01:06.77" resultid="8565" heatid="10778" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="331" swimtime="00:01:22.52" resultid="8566" heatid="10816" lane="0" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="267" swimtime="00:02:38.30" resultid="8567" heatid="10860" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:16.99" />
                    <SPLIT distance="150" swimtime="00:01:57.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="418" swimtime="00:00:35.33" resultid="8568" heatid="10920" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-02" firstname="Mateusz" gender="M" lastname="Stanicki" nation="POL" athleteid="5478">
              <RESULTS>
                <RESULT eventid="1160" points="228" swimtime="00:00:34.19" resultid="8606" heatid="10693" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="1302" points="215" swimtime="00:01:18.20" resultid="8607" heatid="10776" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="187" swimtime="00:02:58.29" resultid="8608" heatid="10859" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="150" swimtime="00:02:09.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="189" swimtime="00:06:23.10" resultid="8609" heatid="10939" lane="9" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                    <SPLIT distance="100" swimtime="00:01:24.15" />
                    <SPLIT distance="150" swimtime="00:02:12.45" />
                    <SPLIT distance="200" swimtime="00:03:01.71" />
                    <SPLIT distance="250" swimtime="00:03:52.10" />
                    <SPLIT distance="300" swimtime="00:04:42.90" />
                    <SPLIT distance="350" swimtime="00:05:33.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-20" firstname="Robert" gender="M" lastname="Budek" nation="POL" athleteid="5305">
              <RESULTS>
                <RESULT eventid="1160" points="250" swimtime="00:00:33.18" resultid="8462" heatid="10698" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1242" points="149" swimtime="00:00:45.28" resultid="8463" heatid="10743" lane="2" entrytime="00:00:45.89" />
                <RESULT eventid="1302" points="204" swimtime="00:01:19.61" resultid="8464" heatid="10777" lane="5" entrytime="00:01:13.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" name="Torpedy" number="4">
              <RESULTS>
                <RESULT eventid="1368" points="413" swimtime="00:02:05.39" resultid="8668" heatid="10802" lane="1" entrytime="00:02:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:11.44" />
                    <SPLIT distance="150" swimtime="00:01:40.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5371" number="1" />
                    <RELAYPOSITION athleteid="5509" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5526" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5534" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" name="Motorówki" number="5">
              <RESULTS>
                <RESULT eventid="1368" points="415" swimtime="00:02:05.19" resultid="8669" heatid="10801" lane="5" entrytime="00:02:05.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:04.14" />
                    <SPLIT distance="150" swimtime="00:01:35.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5279" number="1" />
                    <RELAYPOSITION athleteid="5421" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5379" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5467" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" name="Karmazyny" number="6">
              <RESULTS>
                <RESULT eventid="1368" points="427" swimtime="00:02:04.01" resultid="8670" heatid="10802" lane="9" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:03.60" />
                    <SPLIT distance="150" swimtime="00:01:34.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5412" number="1" />
                    <RELAYPOSITION athleteid="5473" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5438" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5492" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" name="Węgorze" number="8">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Mężczyzn w  kat C  160-199  lat" eventid="1518" points="558" swimtime="00:01:43.06" resultid="8672" heatid="10872" lane="3" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.32" />
                    <SPLIT distance="100" swimtime="00:00:52.37" />
                    <SPLIT distance="150" swimtime="00:01:17.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5313" number="1" />
                    <RELAYPOSITION athleteid="5526" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5534" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5396" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" name="Bojki" number="9">
              <RESULTS>
                <RESULT eventid="1518" points="451" swimtime="00:01:50.62" resultid="8673" heatid="10872" lane="1" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.88" />
                    <SPLIT distance="100" swimtime="00:00:53.74" />
                    <SPLIT distance="150" swimtime="00:01:22.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5279" number="1" />
                    <RELAYPOSITION athleteid="5412" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5455" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5473" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" name="Płetwale" number="10">
              <RESULTS>
                <RESULT eventid="1518" points="350" swimtime="00:02:00.32" resultid="8674" heatid="10870" lane="4" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="100" swimtime="00:01:01.75" />
                    <SPLIT distance="150" swimtime="00:01:30.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5438" number="1" />
                    <RELAYPOSITION athleteid="5305" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5426" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5492" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" name="Makrele" number="7">
              <RESULTS>
                <RESULT eventid="1347" points="318" swimtime="00:02:35.67" resultid="8671" heatid="10798" lane="1" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="100" swimtime="00:01:28.50" />
                    <SPLIT distance="150" swimtime="00:02:04.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5546" number="1" />
                    <RELAYPOSITION athleteid="5329" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5518" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5483" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" name="Turboty" number="11">
              <RESULTS>
                <RESULT eventid="1497" points="416" swimtime="00:02:09.22" resultid="8675" heatid="10868" lane="3" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="150" swimtime="00:01:40.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5483" number="1" />
                    <RELAYPOSITION athleteid="5546" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5540" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5515" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" name="Langusty" number="12">
              <RESULTS>
                <RESULT eventid="1497" points="343" swimtime="00:02:17.83" resultid="8676" heatid="10868" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:07.60" />
                    <SPLIT distance="150" swimtime="00:01:44.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5518" number="1" />
                    <RELAYPOSITION athleteid="5522" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5496" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5406" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="Płaszczki" number="1">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  w  kat B  120-159  lat" eventid="1205" swimtime="00:01:50.56" resultid="8665" heatid="10733" lane="5" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.09" />
                    <SPLIT distance="100" swimtime="00:00:53.89" />
                    <SPLIT distance="150" swimtime="00:01:25.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5313" number="1" />
                    <RELAYPOSITION athleteid="5515" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5483" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5534" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="Meduzy" number="2">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:10.81" resultid="8666" heatid="10732" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.33" />
                    <SPLIT distance="150" swimtime="00:01:41.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5462" number="1" />
                    <RELAYPOSITION athleteid="5522" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5496" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5438" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="Pingwiny" number="3">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:21.02" resultid="8667" heatid="10732" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="150" swimtime="00:01:46.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5540" number="1" />
                    <RELAYPOSITION athleteid="5406" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5362" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5305" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" name="Ośniornice" number="12">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:07.57" resultid="8677" heatid="10929" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:03.31" />
                    <SPLIT distance="150" swimtime="00:01:38.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5412" number="1" />
                    <RELAYPOSITION athleteid="5473" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5540" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5515" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="Piotrosze" number="14">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:26.65" resultid="8678" heatid="10928" lane="3" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                    <SPLIT distance="150" swimtime="00:01:50.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5426" number="1" />
                    <RELAYPOSITION athleteid="5421" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5522" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5496" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="Orki" number="15">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:16.56" resultid="8679" heatid="10929" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:13.43" />
                    <SPLIT distance="150" swimtime="00:01:49.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5371" number="1" />
                    <RELAYPOSITION athleteid="5483" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="5546" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5526" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WEZAB" nation="POL" region="SLA" clubid="3526" name="Weteran  Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁODZIMIERZ" street="ŚW.JANA  4A/4" zip="41-803" />
          <ATHLETES>
            <ATHLETE birthdate="1950-05-10" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" license="502611100005" athleteid="3545">
              <RESULTS>
                <RESULT eventid="1144" points="195" swimtime="00:00:40.92" resultid="8771" heatid="10683" lane="8" entrytime="00:00:41.00" />
                <RESULT eventid="1287" points="161" swimtime="00:01:35.66" resultid="8772" heatid="10766" lane="6" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="112" swimtime="00:03:54.19" resultid="8773" heatid="10851" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.84" />
                    <SPLIT distance="100" swimtime="00:01:50.98" />
                    <SPLIT distance="150" swimtime="00:02:55.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1593" points="65" swimtime="00:05:08.47" resultid="8774" heatid="10894" lane="6" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.19" />
                    <SPLIT distance="100" swimtime="00:02:31.80" />
                    <SPLIT distance="150" swimtime="00:03:54.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="502611100009" athleteid="3565">
              <RESULTS>
                <RESULT eventid="1059" points="446" swimtime="00:10:34.30" resultid="8788" heatid="10667" lane="4" entrytime="00:10:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                    <SPLIT distance="150" swimtime="00:01:56.18" />
                    <SPLIT distance="250" swimtime="00:03:16.60" />
                    <SPLIT distance="350" swimtime="00:04:36.43" />
                    <SPLIT distance="450" swimtime="00:05:56.48" />
                    <SPLIT distance="550" swimtime="00:07:16.20" />
                    <SPLIT distance="650" swimtime="00:08:36.53" />
                    <SPLIT distance="750" swimtime="00:09:56.25" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat E  45-49  lat" eventid="1257" points="416" swimtime="00:03:06.34" resultid="8789" heatid="10756" lane="1" entrytime="00:03:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:30.14" />
                    <SPLIT distance="150" swimtime="00:02:17.58" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters  Kobiet w  kat E  45-49  lat" eventid="1376" points="416" swimtime="00:01:26.18" resultid="8790" heatid="10808" lane="2" entrytime="00:01:24.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat E  45-49  lat" eventid="1525" points="439" swimtime="00:05:50.44" resultid="8791" heatid="10875" lane="2" entrytime="00:05:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:18.60" />
                    <SPLIT distance="150" swimtime="00:02:06.94" />
                    <SPLIT distance="200" swimtime="00:02:54.82" />
                    <SPLIT distance="250" swimtime="00:03:43.88" />
                    <SPLIT distance="300" swimtime="00:04:32.22" />
                    <SPLIT distance="350" swimtime="00:05:12.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="398" swimtime="00:00:40.05" resultid="8792" heatid="10910" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1674" status="DNS" swimtime="00:00:00.00" resultid="8793" heatid="10934" lane="7" entrytime="00:05:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="502611200005" athleteid="8784">
              <RESULTS>
                <RESULT eventid="1160" points="125" swimtime="00:00:41.78" resultid="8785" heatid="10693" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1242" points="72" swimtime="00:00:57.68" resultid="8786" heatid="10743" lane="1" entrytime="00:00:47.50" />
                <RESULT eventid="1422" points="75" swimtime="00:00:53.11" resultid="8787" heatid="10827" lane="5" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="Bastek" nation="POL" license="502611100001" athleteid="3541">
              <RESULTS>
                <RESULT eventid="1144" points="247" swimtime="00:00:37.82" resultid="8768" heatid="10683" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1287" points="207" swimtime="00:01:27.87" resultid="8769" heatid="10767" lane="8" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1674" points="162" swimtime="00:07:12.94" resultid="8770" heatid="10931" lane="5" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                    <SPLIT distance="100" swimtime="00:01:39.50" />
                    <SPLIT distance="150" swimtime="00:02:34.41" />
                    <SPLIT distance="200" swimtime="00:03:30.86" />
                    <SPLIT distance="250" swimtime="00:04:25.77" />
                    <SPLIT distance="300" swimtime="00:05:22.71" />
                    <SPLIT distance="350" swimtime="00:06:18.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-07-16" firstname="Ewald" gender="M" lastname="Bastek" nation="POL" license="502611200001" athleteid="3537">
              <RESULTS>
                <RESULT eventid="1302" points="153" swimtime="00:01:27.53" resultid="8765" heatid="10774" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1482" points="110" swimtime="00:03:32.55" resultid="8766" heatid="10858" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                    <SPLIT distance="100" swimtime="00:01:44.05" />
                    <SPLIT distance="150" swimtime="00:02:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1695" points="133" swimtime="00:07:10.71" resultid="8767" heatid="10937" lane="5" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.80" />
                    <SPLIT distance="100" swimtime="00:01:40.75" />
                    <SPLIT distance="150" swimtime="00:02:36.39" />
                    <SPLIT distance="200" swimtime="00:03:32.75" />
                    <SPLIT distance="250" swimtime="00:04:27.43" />
                    <SPLIT distance="300" swimtime="00:05:24.22" />
                    <SPLIT distance="350" swimtime="00:06:19.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" license="502611100002" athleteid="3531">
              <RESULTS>
                <RESULT eventid="1257" points="171" swimtime="00:04:10.41" resultid="8760" heatid="10753" lane="6" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.09" />
                    <SPLIT distance="100" swimtime="00:02:01.08" />
                    <SPLIT distance="150" swimtime="00:03:07.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="179" swimtime="00:01:54.06" resultid="8761" heatid="10804" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.47" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters Kobiet w  kat J  70-74  lat" eventid="1525" points="102" swimtime="00:09:29.11" resultid="8762" heatid="10873" lane="2" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.94" />
                    <SPLIT distance="100" swimtime="00:02:17.26" />
                    <SPLIT distance="150" swimtime="00:03:35.65" />
                    <SPLIT distance="200" swimtime="00:04:54.72" />
                    <SPLIT distance="250" swimtime="00:06:03.99" />
                    <SPLIT distance="300" swimtime="00:07:14.31" />
                    <SPLIT distance="350" swimtime="00:08:24.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1562" points="113" swimtime="00:01:54.55" resultid="8763" heatid="10883" lane="8" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="177" swimtime="00:00:52.46" resultid="8764" heatid="10907" lane="9" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-07-27" firstname="Danuta" gender="F" lastname="Skorupa" nation="POL" license="502611100012" athleteid="3555">
              <RESULTS>
                <RESULT eventid="1226" points="56" swimtime="00:01:10.39" resultid="8779" heatid="10734" lane="5" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" license="502611200004" athleteid="3572">
              <RESULTS>
                <RESULT eventid="1242" points="161" swimtime="00:00:44.11" resultid="8794" heatid="10743" lane="4" entrytime="00:00:43.26" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="8795" heatid="10774" lane="6" entrytime="00:01:28.82" />
                <RESULT eventid="1452" points="133" swimtime="00:01:41.40" resultid="8796" heatid="10845" lane="1" entrytime="00:01:39.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="115" swimtime="00:03:49.95" resultid="8797" heatid="10900" lane="2" entrytime="00:03:38.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.09" />
                    <SPLIT distance="100" swimtime="00:01:50.21" />
                    <SPLIT distance="150" swimtime="00:02:50.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="Barucha" nation="POL" license="502611200008" athleteid="3550">
              <RESULTS>
                <RESULT eventid="1160" points="276" swimtime="00:00:32.10" resultid="8775" heatid="10698" lane="3" entrytime="00:00:31.68" />
                <RESULT eventid="1242" points="181" swimtime="00:00:42.49" resultid="8776" heatid="10745" lane="0" entrytime="00:00:40.24" />
                <RESULT eventid="1452" points="184" swimtime="00:01:31.07" resultid="8777" heatid="10846" lane="6" entrytime="00:01:28.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="165" swimtime="00:03:23.72" resultid="8778" heatid="10901" lane="2" entrytime="00:03:15.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                    <SPLIT distance="100" swimtime="00:01:40.08" />
                    <SPLIT distance="150" swimtime="00:02:32.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" license="502611200002" athleteid="3527">
              <RESULTS>
                <RESULT eventid="1272" points="188" swimtime="00:03:41.56" resultid="8757" heatid="10758" lane="4" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.70" />
                    <SPLIT distance="100" swimtime="00:01:48.93" />
                    <SPLIT distance="150" swimtime="00:02:47.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="177" swimtime="00:01:41.67" resultid="8758" heatid="10811" lane="6" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="193" swimtime="00:00:45.70" resultid="8759" heatid="10915" lane="8" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-28" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="502611200007" athleteid="8780">
              <RESULTS>
                <RESULT eventid="1160" points="208" swimtime="00:00:35.24" resultid="8781" heatid="10697" lane="3" entrytime="00:00:32.56" />
                <RESULT eventid="1302" points="189" swimtime="00:01:21.64" resultid="8782" heatid="10777" lane="7" entrytime="00:01:15.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="224" swimtime="00:00:36.92" resultid="8783" heatid="10829" lane="8" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1368" points="173" swimtime="00:02:47.60" resultid="8801" heatid="10800" lane="1" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="150" swimtime="00:01:03.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3550" number="1" />
                    <RELAYPOSITION athleteid="3527" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="8780" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3537" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1518" points="164" swimtime="00:02:34.77" resultid="8803" heatid="10870" lane="8" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="150" swimtime="00:01:59.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3527" number="1" />
                    <RELAYPOSITION athleteid="8784" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3572" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="8780" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1347" points="218" swimtime="00:02:56.66" resultid="8800" heatid="10798" lane="8" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.42" />
                    <SPLIT distance="100" swimtime="00:01:40.81" />
                    <SPLIT distance="150" swimtime="00:02:15.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3541" number="1" />
                    <RELAYPOSITION athleteid="3531" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3565" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3545" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="5">
              <RESULTS>
                <RESULT eventid="1497" points="203" swimtime="00:02:44.20" resultid="8802" heatid="10868" lane="5" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:29.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3541" number="1" />
                    <RELAYPOSITION athleteid="3531" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3545" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3565" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:43.77" resultid="8798" heatid="10731" lane="5" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                    <SPLIT distance="100" swimtime="00:01:27.98" />
                    <SPLIT distance="150" swimtime="00:02:09.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3541" number="1" />
                    <RELAYPOSITION athleteid="3531" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="8784" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="8780" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1205" swimtime="00:02:23.47" resultid="8799" heatid="10732" lane="0" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:01:19.09" />
                    <SPLIT distance="150" swimtime="00:01:51.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3545" number="1" />
                    <RELAYPOSITION athleteid="3537" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3565" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3550" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:55.53" resultid="8804" heatid="10927" lane="4" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                    <SPLIT distance="100" swimtime="00:01:39.88" />
                    <SPLIT distance="150" swimtime="00:02:16.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3572" number="1" />
                    <RELAYPOSITION athleteid="3531" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="8780" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3541" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="8">
              <RESULTS>
                <RESULT eventid="1653" swimtime="00:02:45.58" resultid="8805" heatid="10928" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:02.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3550" number="1" />
                    <RELAYPOSITION athleteid="3527" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3565" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3545" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WSBDG" nation="POL" region="11" clubid="10613" name="WSB Dąbrowa Górnicza">
          <ATHLETES>
            <ATHLETE birthdate="1993-01-01" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" athleteid="10111">
              <RESULTS>
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="10112" heatid="10672" lane="9" entrytime="00:11:20.00" />
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="10113" heatid="10703" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="10114" heatid="10723" lane="6" entrytime="00:03:00.00" />
                <RESULT eventid="1242" points="282" swimtime="00:00:36.64" resultid="10115" heatid="10750" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1272" points="241" swimtime="00:03:23.94" resultid="10116" heatid="10762" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                    <SPLIT distance="100" swimtime="00:01:35.02" />
                    <SPLIT distance="150" swimtime="00:02:28.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="313" swimtime="00:01:24.12" resultid="10117" heatid="10816" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" status="DNS" swimtime="00:00:00.00" resultid="10118" heatid="10849" lane="6" entrytime="00:01:08.00" />
                <RESULT eventid="1608" points="227" swimtime="00:03:03.33" resultid="10119" heatid="10902" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                    <SPLIT distance="100" swimtime="00:01:27.29" />
                    <SPLIT distance="150" swimtime="00:02:14.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="430" swimtime="00:00:34.99" resultid="10120" heatid="10925" lane="3" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WSHS" nation="POL" region="11" clubid="10614" name="Wyższa Szkoła Humanitas Sosnowiec">
          <ATHLETES>
            <ATHLETE birthdate="1996-01-01" firstname="Kinga" gender="F" lastname="Pluta" nation="POL" athleteid="10121">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="10122" heatid="10667" lane="7" entrytime="00:12:30.00" />
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="10123" heatid="10687" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="10124" heatid="10715" lane="2" entrytime="00:03:15.00" />
                <RESULT eventid="1226" points="359" swimtime="00:00:38.05" resultid="10125" heatid="10739" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1257" points="363" swimtime="00:03:14.84" resultid="10126" heatid="10755" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.14" />
                    <SPLIT distance="100" swimtime="00:01:32.98" />
                    <SPLIT distance="150" swimtime="00:02:24.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="413" swimtime="00:01:26.39" resultid="10127" heatid="10807" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="10128" heatid="10841" lane="0" entrytime="00:01:30.00" />
                <RESULT eventid="1593" points="335" swimtime="00:02:58.47" resultid="10129" heatid="10896" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                    <SPLIT distance="100" swimtime="00:01:28.23" />
                    <SPLIT distance="150" swimtime="00:02:13.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1623" points="450" swimtime="00:00:38.45" resultid="10130" heatid="10911" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ZKDRZ" nation="POL" region="LBS" clubid="4058" name="ZKS Drzonków">
          <CONTACT email="llfpiotr@gmail.com" name="Barta Piotr" phone="602347348" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-18" firstname="Piotr" gender="M" lastname="Barta" nation="POL" athleteid="4059">
              <RESULTS>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="6420" heatid="10729" lane="0" entrytime="00:02:32.00" entrycourse="LCM" />
                <RESULT eventid="1272" points="491" swimtime="00:02:40.98" resultid="6421" heatid="10764" lane="2" entrytime="00:02:38.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:01:16.80" />
                    <SPLIT distance="150" swimtime="00:01:58.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="467" swimtime="00:01:13.62" resultid="6422" heatid="10818" lane="5" entrytime="00:01:13.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="6424" heatid="10924" lane="4" entrytime="00:00:33.33" entrycourse="LCM" />
                <RESULT eventid="1695" status="DNS" swimtime="00:00:00.00" resultid="6425" heatid="10944" lane="3" entrytime="00:04:47.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ZUBR" nation="BLR" clubid="3607" name="Zubr">
          <CONTACT email="pr3429@gmail.com" name="Minsk Masters Swimming Club ZUBR" phone="+375445313201" />
          <ATHLETES>
            <ATHLETE birthdate="1972-01-02" firstname="Aliaksandr" gender="M" lastname="Puzan" nation="BLR" athleteid="3814">
              <RESULTS>
                <RESULT eventid="1160" points="435" swimtime="00:00:27.59" resultid="10167" heatid="10704" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="1302" points="423" swimtime="00:01:02.46" resultid="10168" heatid="10785" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="371" swimtime="00:00:31.20" resultid="10169" heatid="10833" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="1578" points="338" swimtime="00:01:11.47" resultid="10170" heatid="10889" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-12" firstname="Roman12021974" gender="M" lastname="Kostitsin" nation="BLR" athleteid="9039">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="10157" heatid="10700" lane="5" entrytime="00:00:30.10" entrycourse="LCM" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="10158" heatid="10761" lane="4" entrytime="00:03:02.17" entrycourse="LCM" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="10159" heatid="10816" lane="9" entrytime="00:01:22.60" entrycourse="LCM" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="10160" heatid="10830" lane="1" entrytime="00:00:34.15" entrycourse="LCM" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="10161" heatid="10922" lane="0" entrytime="00:00:36.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-05-10" firstname="Siarhei" gender="M" lastname="Aliashkevich" nation="BLR" athleteid="9045">
              <RESULTS>
                <RESULT eventid="1190" points="419" swimtime="00:02:32.31" resultid="10162" heatid="10728" lane="6" entrytime="00:02:34.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:10.87" />
                    <SPLIT distance="150" swimtime="00:01:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="449" swimtime="00:00:31.38" resultid="10163" heatid="10749" lane="5" entrytime="00:00:31.66" entrycourse="LCM" />
                <RESULT eventid="1422" points="408" swimtime="00:00:30.22" resultid="10164" heatid="10835" lane="8" entrytime="00:00:29.67" entrycourse="LCM" />
                <RESULT eventid="1452" points="397" swimtime="00:01:10.50" resultid="10165" heatid="10849" lane="1" entrytime="00:01:09.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="392" swimtime="00:02:32.86" resultid="10166" heatid="10904" lane="9" entrytime="00:02:34.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                    <SPLIT distance="100" swimtime="00:01:14.57" />
                    <SPLIT distance="150" swimtime="00:01:54.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SKPPR" nation="SVK" region="VSO" clubid="2949" name="Športový klub polície Prešov">
          <CONTACT city="Prešov" email="jzpl@centrum.sk" name="Žilinský Jozef" state="SVK" street="Mirka Nešpora 17" zip="080 01" />
          <ATHLETES>
            <ATHLETE birthdate="1952-03-23" firstname="Jozef" gender="M" lastname="Žilinský" nation="SVK" license="SVK11472" athleteid="2950">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="7911" heatid="10691" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1242" status="DNS" swimtime="00:00:00.00" resultid="7912" heatid="10742" lane="8" entrytime="00:00:54.25" />
                <RESULT eventid="1392" status="DNS" swimtime="00:00:00.00" resultid="7913" heatid="10810" lane="7" entrytime="00:01:58.57" />
                <RESULT eventid="1452" status="DNS" swimtime="00:00:00.00" resultid="7914" heatid="10844" lane="2" entrytime="00:02:09.57" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="7915" heatid="10914" lane="0" entrytime="00:00:50.31" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="MTP Delfin Cieszyn" version="Build 22680">
    <CONTACT name="GeoLogix AG" street="Muristrasse 60" city="Bern" zip="3006" country="CH" phone="+41 31 356 80 56" fax="+41 31 356 80 81" email="info@splash-software.ch" internet="http://www.splash-software.ch" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Katowice" name="Zimowe Otwarte Mistrzostwa Polski Masters" course="SCM" deadline="2012-11-14" hostclub="UKS Wodnik 29 Katowice" hostclub.url="http://www.wodnik29.pl" nation="POL" organizer="UKS Wodnik 29 Katowice" organizer.url="http://www.wodnik29.pl" timing="AUTOMATIC">
      <AGEDATE value="2012-11-23" type="YEAR" />
      <POOL lanemin="1" lanemax="6" />
      <POINTTABLE pointtableid="1008" name="DSV Master Performance Table" version="2004" />
      <CONTACT city="Katowice" email="kontakt@delfincieszyn.pl" name="Łukasz Widzik" phone="660749175" street="Mikołowska 72" />
      <SESSIONS>
        <SESSION date="2012-11-23" daytime="16:00" name="Blok I" number="1" warmupfrom="15:00">
          <EVENTS>
            <EVENT eventid="1058" daytime="16:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1060" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1061" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4038" />
                    <RANKING order="2" place="2" resultid="4418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2034" />
                    <RANKING order="2" place="2" resultid="2387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2790" />
                    <RANKING order="2" place="2" resultid="4046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4194" />
                    <RANKING order="2" place="2" resultid="2291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3799" />
                    <RANKING order="2" place="2" resultid="2558" />
                    <RANKING order="3" place="3" resultid="2787" />
                    <RANKING order="4" place="-1" resultid="4791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3835" />
                    <RANKING order="2" place="2" resultid="3776" />
                    <RANKING order="3" place="3" resultid="1988" />
                    <RANKING order="4" place="-1" resultid="1957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="69" agemin="65" name="I: 65 - 69 lat" />
                <AGEGROUP agegroupid="1070" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1071" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1072" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1073" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6428" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6429" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6430" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6431" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="16:30" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2016" />
                    <RANKING order="2" place="2" resultid="4611" />
                    <RANKING order="3" place="3" resultid="4003" />
                    <RANKING order="4" place="-1" resultid="1732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2422" />
                    <RANKING order="2" place="2" resultid="2455" />
                    <RANKING order="3" place="3" resultid="4763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4706" />
                    <RANKING order="2" place="2" resultid="2504" />
                    <RANKING order="3" place="3" resultid="3372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1096" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2489" />
                    <RANKING order="2" place="2" resultid="2574" />
                    <RANKING order="3" place="3" resultid="4812" />
                    <RANKING order="4" place="4" resultid="3179" />
                    <RANKING order="5" place="5" resultid="2550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4001" />
                    <RANKING order="2" place="2" resultid="3448" />
                    <RANKING order="3" place="3" resultid="2520" />
                    <RANKING order="4" place="4" resultid="1741" />
                    <RANKING order="5" place="5" resultid="3228" />
                    <RANKING order="6" place="6" resultid="3119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3545" />
                    <RANKING order="2" place="2" resultid="2680" />
                    <RANKING order="3" place="3" resultid="2379" />
                    <RANKING order="4" place="4" resultid="3538" />
                    <RANKING order="5" place="5" resultid="2566" />
                    <RANKING order="6" place="6" resultid="2402" />
                    <RANKING order="7" place="7" resultid="3250" />
                    <RANKING order="8" place="8" resultid="1869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4800" />
                    <RANKING order="2" place="2" resultid="2528" />
                    <RANKING order="3" place="3" resultid="3039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2712" />
                    <RANKING order="2" place="2" resultid="3961" />
                    <RANKING order="3" place="3" resultid="2916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4586" />
                    <RANKING order="2" place="2" resultid="2512" />
                    <RANKING order="3" place="3" resultid="1951" />
                    <RANKING order="4" place="4" resultid="3212" />
                    <RANKING order="5" place="5" resultid="3909" />
                    <RANKING order="6" place="6" resultid="3812" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2634" />
                    <RANKING order="2" place="2" resultid="3947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3204" />
                    <RANKING order="2" place="2" resultid="3852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4290" />
                    <RANKING order="2" place="2" resultid="3696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6485" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6486" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6487" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6488" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6489" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6490" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6491" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6492" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="17:40" gender="X" number="3" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2318" />
                    <RANKING order="2" place="2" resultid="3499" />
                    <RANKING order="3" place="3" resultid="4123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2320" />
                    <RANKING order="2" place="2" resultid="2795" />
                    <RANKING order="3" place="3" resultid="4125" />
                    <RANKING order="4" place="4" resultid="4483" />
                    <RANKING order="5" place="5" resultid="4484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1942" />
                    <RANKING order="2" place="2" resultid="2319" />
                    <RANKING order="3" place="3" resultid="3986" />
                    <RANKING order="4" place="4" resultid="4250" />
                    <RANKING order="5" place="5" resultid="2322" />
                    <RANKING order="6" place="6" resultid="3163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2005" />
                    <RANKING order="2" place="2" resultid="4249" />
                    <RANKING order="3" place="3" resultid="2321" />
                    <RANKING order="4" place="-1" resultid="1889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="-1" agemin="280" name="F: 280 lat i starsi" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6494" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6495" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6496" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6497" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1122" daytime="17:55" gender="F" number="4" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1123" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2025" />
                    <RANKING order="2" place="2" resultid="6029" />
                    <RANKING order="3" place="3" resultid="3624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4570" />
                    <RANKING order="2" place="2" resultid="2698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4054" />
                    <RANKING order="2" place="2" resultid="3477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1657" />
                    <RANKING order="2" place="2" resultid="2791" />
                    <RANKING order="3" place="3" resultid="2146" />
                    <RANKING order="4" place="4" resultid="3045" />
                    <RANKING order="5" place="-1" resultid="4298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4411" />
                    <RANKING order="2" place="2" resultid="4226" />
                    <RANKING order="3" place="3" resultid="4110" />
                    <RANKING order="4" place="4" resultid="3294" />
                    <RANKING order="5" place="5" resultid="2879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4792" />
                    <RANKING order="2" place="2" resultid="2409" />
                    <RANKING order="3" place="3" resultid="4578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1944" />
                    <RANKING order="2" place="2" resultid="3141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2952" />
                    <RANKING order="2" place="2" resultid="4437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1132" agemax="69" agemin="65" name="I: 65 - 69 lat" />
                <AGEGROUP agegroupid="1133" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1134" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1135" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6441" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6442" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6443" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6444" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6445" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1137" daytime="19:15" gender="M" number="5" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1138" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4703" />
                    <RANKING order="2" place="2" resultid="3873" />
                    <RANKING order="3" place="3" resultid="4561" />
                    <RANKING order="4" place="4" resultid="2073" />
                    <RANKING order="5" place="5" resultid="4550" />
                    <RANKING order="6" place="-1" resultid="4594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4632" />
                    <RANKING order="2" place="2" resultid="3882" />
                    <RANKING order="3" place="3" resultid="6498" />
                    <RANKING order="4" place="4" resultid="2081" />
                    <RANKING order="5" place="5" resultid="6500" />
                    <RANKING order="6" place="6" resultid="3410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1140" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3282" />
                    <RANKING order="2" place="2" resultid="3638" />
                    <RANKING order="3" place="3" resultid="3820" />
                    <RANKING order="4" place="4" resultid="4353" />
                    <RANKING order="5" place="5" resultid="2186" />
                    <RANKING order="6" place="-1" resultid="3328" />
                    <RANKING order="7" place="-1" resultid="3336" />
                    <RANKING order="8" place="-1" resultid="1780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1141" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2463" />
                    <RANKING order="2" place="2" resultid="3303" />
                    <RANKING order="3" place="3" resultid="2256" />
                    <RANKING order="4" place="4" resultid="2542" />
                    <RANKING order="5" place="5" resultid="3382" />
                    <RANKING order="6" place="6" resultid="2497" />
                    <RANKING order="7" place="-1" resultid="2894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3167" />
                    <RANKING order="2" place="2" resultid="2474" />
                    <RANKING order="3" place="3" resultid="3826" />
                    <RANKING order="4" place="4" resultid="6038" />
                    <RANKING order="5" place="5" resultid="2042" />
                    <RANKING order="6" place="6" resultid="3865" />
                    <RANKING order="7" place="7" resultid="3242" />
                    <RANKING order="8" place="8" resultid="4323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4374" />
                    <RANKING order="2" place="2" resultid="4656" />
                    <RANKING order="3" place="3" resultid="2270" />
                    <RANKING order="4" place="4" resultid="2282" />
                    <RANKING order="5" place="-1" resultid="2692" />
                    <RANKING order="6" place="-1" resultid="2167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4005" />
                    <RANKING order="2" place="2" resultid="1800" />
                    <RANKING order="3" place="3" resultid="3319" />
                    <RANKING order="4" place="4" resultid="2175" />
                    <RANKING order="5" place="5" resultid="4403" />
                    <RANKING order="6" place="-1" resultid="2064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2759" />
                    <RANKING order="2" place="2" resultid="3844" />
                    <RANKING order="3" place="3" resultid="2764" />
                    <RANKING order="4" place="4" resultid="4140" />
                    <RANKING order="5" place="5" resultid="3220" />
                    <RANKING order="6" place="6" resultid="6039" />
                    <RANKING order="7" place="7" resultid="3053" />
                    <RANKING order="8" place="8" resultid="3149" />
                    <RANKING order="9" place="-1" resultid="3184" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4471" />
                    <RANKING order="2" place="2" resultid="2121" />
                    <RANKING order="3" place="3" resultid="3955" />
                    <RANKING order="4" place="4" resultid="2980" />
                    <RANKING order="5" place="5" resultid="2618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2230" />
                    <RANKING order="2" place="2" resultid="4366" />
                    <RANKING order="3" place="3" resultid="2986" />
                    <RANKING order="4" place="-1" resultid="2197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1149" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1662" />
                    <RANKING order="2" place="2" resultid="2623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6514" agemax="89" agemin="85" name="M: 85 - 89 lat" />
                <AGEGROUP agegroupid="1151" agemax="-1" agemin="90" name="N: 90 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1863" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6446" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6447" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6448" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6449" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6450" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6451" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6452" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6453" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6454" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6455" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6456" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6457" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2012-11-24" daytime="09:00" name="Blok II" number="2" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1153" daytime="09:00" gender="F" number="6" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1154" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2098" />
                    <RANKING order="2" place="2" resultid="2447" />
                    <RANKING order="3" place="3" resultid="3625" />
                    <RANKING order="4" place="4" resultid="2721" />
                    <RANKING order="5" place="-1" resultid="2646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3310" />
                    <RANKING order="2" place="2" resultid="2277" />
                    <RANKING order="3" place="3" resultid="4085" />
                    <RANKING order="4" place="4" resultid="4571" />
                    <RANKING order="5" place="5" resultid="4419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2856" />
                    <RANKING order="2" place="2" resultid="4683" />
                    <RANKING order="3" place="3" resultid="3632" />
                    <RANKING order="4" place="4" resultid="2035" />
                    <RANKING order="5" place="5" resultid="4597" />
                    <RANKING order="6" place="6" resultid="2388" />
                    <RANKING order="7" place="7" resultid="4447" />
                    <RANKING order="8" place="8" resultid="4055" />
                    <RANKING order="9" place="9" resultid="3512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3610" />
                    <RANKING order="2" place="2" resultid="3524" />
                    <RANKING order="3" place="3" resultid="3995" />
                    <RANKING order="4" place="-1" resultid="2147" />
                    <RANKING order="5" place="-1" resultid="2839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4479" />
                    <RANKING order="2" place="2" resultid="4208" />
                    <RANKING order="3" place="3" resultid="2292" />
                    <RANKING order="4" place="-1" resultid="4111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2130" />
                    <RANKING order="2" place="2" resultid="4664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1844" />
                    <RANKING order="2" place="2" resultid="1838" />
                    <RANKING order="3" place="3" resultid="3836" />
                    <RANKING order="4" place="4" resultid="3777" />
                    <RANKING order="5" place="5" resultid="1999" />
                    <RANKING order="6" place="6" resultid="3617" />
                    <RANKING order="7" place="7" resultid="3471" />
                    <RANKING order="8" place="8" resultid="1989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2219" />
                    <RANKING order="2" place="2" resultid="1821" />
                    <RANKING order="3" place="3" resultid="1972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4165" />
                    <RANKING order="2" place="2" resultid="1875" />
                    <RANKING order="3" place="3" resultid="2154" />
                    <RANKING order="4" place="4" resultid="1965" />
                    <RANKING order="5" place="5" resultid="2953" />
                    <RANKING order="6" place="6" resultid="4189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4220" />
                    <RANKING order="2" place="2" resultid="2160" />
                    <RANKING order="3" place="3" resultid="2960" />
                    <RANKING order="4" place="-1" resultid="4457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4640" />
                    <RANKING order="2" place="2" resultid="1813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1166" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1167" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6074" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6075" daytime="09:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6076" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6077" daytime="09:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6078" daytime="09:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6079" daytime="09:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6080" daytime="09:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6081" daytime="09:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6082" daytime="09:20" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1168" daytime="09:20" gender="M" number="7" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1169" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3874" />
                    <RANKING order="2" place="2" resultid="2799" />
                    <RANKING order="3" place="3" resultid="4612" />
                    <RANKING order="4" place="4" resultid="2017" />
                    <RANKING order="5" place="5" resultid="2212" />
                    <RANKING order="6" place="6" resultid="4529" />
                    <RANKING order="7" place="-1" resultid="3062" />
                    <RANKING order="8" place="-1" resultid="4544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3100" />
                    <RANKING order="2" place="2" resultid="3108" />
                    <RANKING order="3" place="3" resultid="4554" />
                    <RANKING order="4" place="4" resultid="2725" />
                    <RANKING order="5" place="5" resultid="3396" />
                    <RANKING order="6" place="6" resultid="4312" />
                    <RANKING order="7" place="7" resultid="2651" />
                    <RANKING order="8" place="8" resultid="1793" />
                    <RANKING order="9" place="9" resultid="2662" />
                    <RANKING order="10" place="10" resultid="3460" />
                    <RANKING order="11" place="11" resultid="3785" />
                    <RANKING order="12" place="12" resultid="3411" />
                    <RANKING order="13" place="13" resultid="2582" />
                    <RANKING order="14" place="14" resultid="4104" />
                    <RANKING order="15" place="-1" resultid="2666" />
                    <RANKING order="16" place="-1" resultid="2733" />
                    <RANKING order="17" place="-1" resultid="3070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4443" />
                    <RANKING order="2" place="2" resultid="3639" />
                    <RANKING order="3" place="3" resultid="4707" />
                    <RANKING order="4" place="4" resultid="1781" />
                    <RANKING order="5" place="5" resultid="3329" />
                    <RANKING order="6" place="6" resultid="4244" />
                    <RANKING order="7" place="7" resultid="4073" />
                    <RANKING order="8" place="8" resultid="3361" />
                    <RANKING order="9" place="9" resultid="4354" />
                    <RANKING order="10" place="10" resultid="3403" />
                    <RANKING order="11" place="-1" resultid="3344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2490" />
                    <RANKING order="2" place="2" resultid="2575" />
                    <RANKING order="3" place="3" resultid="4023" />
                    <RANKING order="4" place="4" resultid="4813" />
                    <RANKING order="5" place="5" resultid="3383" />
                    <RANKING order="6" place="6" resultid="2848" />
                    <RANKING order="7" place="7" resultid="2551" />
                    <RANKING order="8" place="8" resultid="3456" />
                    <RANKING order="9" place="9" resultid="2396" />
                    <RANKING order="10" place="10" resultid="4604" />
                    <RANKING order="11" place="-1" resultid="2895" />
                    <RANKING order="12" place="-1" resultid="3980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2049" />
                    <RANKING order="2" place="2" resultid="1750" />
                    <RANKING order="3" place="3" resultid="2475" />
                    <RANKING order="4" place="4" resultid="2521" />
                    <RANKING order="5" place="5" resultid="1996" />
                    <RANKING order="6" place="6" resultid="3120" />
                    <RANKING order="7" place="7" resultid="3229" />
                    <RANKING order="8" place="8" resultid="2441" />
                    <RANKING order="9" place="9" resultid="3974" />
                    <RANKING order="10" place="10" resultid="4324" />
                    <RANKING order="11" place="-1" resultid="3891" />
                    <RANKING order="12" place="-1" resultid="2843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3546" />
                    <RANKING order="2" place="2" resultid="4331" />
                    <RANKING order="3" place="3" resultid="1936" />
                    <RANKING order="4" place="4" resultid="4080" />
                    <RANKING order="5" place="5" resultid="3251" />
                    <RANKING order="6" place="6" resultid="2168" />
                    <RANKING order="7" place="7" resultid="2283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4031" />
                    <RANKING order="2" place="2" resultid="4305" />
                    <RANKING order="3" place="3" resultid="4801" />
                    <RANKING order="4" place="4" resultid="3495" />
                    <RANKING order="5" place="5" resultid="2245" />
                    <RANKING order="6" place="6" resultid="6032" />
                    <RANKING order="7" place="7" resultid="3040" />
                    <RANKING order="8" place="8" resultid="4404" />
                    <RANKING order="9" place="-1" resultid="1801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4360" />
                    <RANKING order="2" place="2" resultid="2743" />
                    <RANKING order="3" place="3" resultid="3768" />
                    <RANKING order="4" place="4" resultid="3659" />
                    <RANKING order="5" place="5" resultid="3704" />
                    <RANKING order="6" place="6" resultid="4141" />
                    <RANKING order="7" place="7" resultid="3962" />
                    <RANKING order="8" place="8" resultid="3734" />
                    <RANKING order="9" place="9" resultid="2057" />
                    <RANKING order="10" place="10" resultid="3221" />
                    <RANKING order="11" place="11" resultid="3001" />
                    <RANKING order="12" place="12" resultid="2906" />
                    <RANKING order="13" place="13" resultid="3150" />
                    <RANKING order="14" place="-1" resultid="3531" />
                    <RANKING order="15" place="-1" resultid="4066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4587" />
                    <RANKING order="2" place="2" resultid="3583" />
                    <RANKING order="3" place="3" resultid="2513" />
                    <RANKING order="4" place="4" resultid="3813" />
                    <RANKING order="5" place="5" resultid="4215" />
                    <RANKING order="6" place="6" resultid="3910" />
                    <RANKING order="7" place="7" resultid="3008" />
                    <RANKING order="8" place="-1" resultid="2981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2635" />
                    <RANKING order="2" place="2" resultid="3948" />
                    <RANKING order="3" place="3" resultid="3941" />
                    <RANKING order="4" place="4" resultid="2204" />
                    <RANKING order="5" place="5" resultid="2987" />
                    <RANKING order="6" place="-1" resultid="2198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6083" daytime="09:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6084" daytime="09:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6085" daytime="09:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6086" daytime="09:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6087" daytime="09:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6088" daytime="09:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6089" daytime="09:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6090" daytime="09:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6091" daytime="09:40" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6092" daytime="09:40" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6093" daytime="09:40" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6094" daytime="09:45" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6095" daytime="09:45" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6096" daytime="09:45" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="6097" daytime="09:50" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="6098" daytime="09:50" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="6099" daytime="09:50" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="6100" daytime="09:55" number="18" order="18" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" daytime="09:55" gender="F" number="8" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1184" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2099" />
                    <RANKING order="2" place="2" resultid="4778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3652" />
                    <RANKING order="2" place="2" resultid="4425" />
                    <RANKING order="3" place="3" resultid="2208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3611" />
                    <RANKING order="2" place="2" resultid="3265" />
                    <RANKING order="3" place="3" resultid="3046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4195" />
                    <RANKING order="2" place="2" resultid="3258" />
                    <RANKING order="3" place="3" resultid="3295" />
                    <RANKING order="4" place="4" resultid="2260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4380" />
                    <RANKING order="2" place="2" resultid="4793" />
                    <RANKING order="3" place="3" resultid="2559" />
                    <RANKING order="4" place="4" resultid="4579" />
                    <RANKING order="5" place="5" resultid="4452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2142" />
                    <RANKING order="2" place="2" resultid="4678" />
                    <RANKING order="3" place="3" resultid="1958" />
                    <RANKING order="4" place="4" resultid="3465" />
                    <RANKING order="5" place="5" resultid="3142" />
                    <RANKING order="6" place="6" resultid="2994" />
                    <RANKING order="7" place="-1" resultid="4228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3936" />
                    <RANKING order="2" place="2" resultid="1973" />
                    <RANKING order="3" place="3" resultid="3134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2155" />
                    <RANKING order="2" place="2" resultid="2807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4176" />
                    <RANKING order="2" place="2" resultid="4152" />
                    <RANKING order="3" place="3" resultid="2931" />
                    <RANKING order="4" place="4" resultid="2161" />
                    <RANKING order="5" place="5" resultid="6539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6511" />
                    <RANKING order="2" place="2" resultid="4651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1197" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6101" daytime="09:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6102" daytime="10:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6103" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6104" daytime="10:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6105" daytime="10:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6106" daytime="10:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6107" daytime="10:25" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1198" daytime="10:30" gender="M" number="9" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1199" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4562" />
                    <RANKING order="2" place="2" resultid="4534" />
                    <RANKING order="3" place="3" resultid="3793" />
                    <RANKING order="4" place="-1" resultid="1733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4555" />
                    <RANKING order="2" place="2" resultid="4538" />
                    <RANKING order="3" place="3" resultid="4463" />
                    <RANKING order="4" place="4" resultid="2114" />
                    <RANKING order="5" place="5" resultid="3277" />
                    <RANKING order="6" place="6" resultid="3390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2505" />
                    <RANKING order="2" place="2" resultid="3330" />
                    <RANKING order="3" place="3" resultid="3337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2576" />
                    <RANKING order="2" place="2" resultid="2543" />
                    <RANKING order="3" place="3" resultid="2315" />
                    <RANKING order="4" place="4" resultid="2498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3449" />
                    <RANKING order="2" place="2" resultid="3014" />
                    <RANKING order="3" place="3" resultid="1742" />
                    <RANKING order="4" place="4" resultid="3243" />
                    <RANKING order="5" place="-1" resultid="4011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3505" />
                    <RANKING order="2" place="2" resultid="3968" />
                    <RANKING order="3" place="3" resultid="3539" />
                    <RANKING order="4" place="4" resultid="4338" />
                    <RANKING order="5" place="-1" resultid="2380" />
                    <RANKING order="6" place="-1" resultid="2693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3552" />
                    <RANKING order="2" place="2" resultid="4625" />
                    <RANKING order="3" place="3" resultid="2536" />
                    <RANKING order="4" place="4" resultid="2176" />
                    <RANKING order="5" place="-1" resultid="1881" />
                    <RANKING order="6" place="-1" resultid="3320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2744" />
                    <RANKING order="2" place="2" resultid="2713" />
                    <RANKING order="3" place="3" resultid="1831" />
                    <RANKING order="4" place="4" resultid="3054" />
                    <RANKING order="5" place="5" resultid="3845" />
                    <RANKING order="6" place="6" resultid="2917" />
                    <RANKING order="7" place="7" resultid="3151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4588" />
                    <RANKING order="2" place="2" resultid="1827" />
                    <RANKING order="3" place="3" resultid="2514" />
                    <RANKING order="4" place="4" resultid="1952" />
                    <RANKING order="5" place="5" resultid="3213" />
                    <RANKING order="6" place="6" resultid="3570" />
                    <RANKING order="7" place="7" resultid="2301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3949" />
                    <RANKING order="2" place="2" resultid="2688" />
                    <RANKING order="3" place="3" resultid="2988" />
                    <RANKING order="4" place="4" resultid="2812" />
                    <RANKING order="5" place="-1" resultid="2973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4181" />
                    <RANKING order="2" place="2" resultid="3157" />
                    <RANKING order="3" place="3" resultid="1982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6108" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6109" daytime="10:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6110" daytime="10:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6111" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6112" daytime="10:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6113" daytime="10:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6114" daytime="11:00" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6115" daytime="11:00" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6116" daytime="11:05" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6117" daytime="11:10" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1213" daytime="11:10" gender="F" number="10" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1214" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2705" />
                    <RANKING order="2" place="2" resultid="2448" />
                    <RANKING order="3" place="3" resultid="2026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3311" />
                    <RANKING order="2" place="2" resultid="2238" />
                    <RANKING order="3" place="3" resultid="4039" />
                    <RANKING order="4" place="4" resultid="4690" />
                    <RANKING order="5" place="5" resultid="1921" />
                    <RANKING order="6" place="6" resultid="4019" />
                    <RANKING order="7" place="-1" resultid="2887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3633" />
                    <RANKING order="2" place="2" resultid="2389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4299" />
                    <RANKING order="2" place="2" resultid="4236" />
                    <RANKING order="3" place="3" resultid="3996" />
                    <RANKING order="4" place="4" resultid="4389" />
                    <RANKING order="5" place="5" resultid="4047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4209" />
                    <RANKING order="2" place="2" resultid="4412" />
                    <RANKING order="3" place="3" resultid="2293" />
                    <RANKING order="4" place="4" resultid="4112" />
                    <RANKING order="5" place="5" resultid="3296" />
                    <RANKING order="6" place="6" resultid="2261" />
                    <RANKING order="7" place="7" resultid="2880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2131" />
                    <RANKING order="2" place="2" resultid="2410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1839" />
                    <RANKING order="2" place="2" resultid="3837" />
                    <RANKING order="3" place="3" resultid="1768" />
                    <RANKING order="4" place="4" resultid="1945" />
                    <RANKING order="5" place="5" resultid="3618" />
                    <RANKING order="6" place="6" resultid="2995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4147" />
                    <RANKING order="2" place="2" resultid="3135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4166" />
                    <RANKING order="2" place="2" resultid="2770" />
                    <RANKING order="3" place="3" resultid="2938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4172" />
                    <RANKING order="2" place="2" resultid="4221" />
                    <RANKING order="3" place="3" resultid="2945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4641" />
                    <RANKING order="2" place="2" resultid="1814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6118" daytime="11:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6119" daytime="11:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6120" daytime="11:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6121" daytime="11:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6122" daytime="11:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6123" daytime="11:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6124" daytime="11:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6125" daytime="11:20" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1228" daytime="11:25" gender="M" number="11" order="13" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1229" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2751" />
                    <RANKING order="2" place="2" resultid="2800" />
                    <RANKING order="3" place="3" resultid="2863" />
                    <RANKING order="4" place="4" resultid="4613" />
                    <RANKING order="5" place="5" resultid="2655" />
                    <RANKING order="6" place="6" resultid="4545" />
                    <RANKING order="7" place="7" resultid="2417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3109" />
                    <RANKING order="2" place="2" resultid="2629" />
                    <RANKING order="3" place="3" resultid="4432" />
                    <RANKING order="4" place="4" resultid="3397" />
                    <RANKING order="5" place="5" resultid="3391" />
                    <RANKING order="6" place="-1" resultid="2734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3283" />
                    <RANKING order="2" place="2" resultid="3604" />
                    <RANKING order="3" place="3" resultid="4708" />
                    <RANKING order="4" place="4" resultid="2089" />
                    <RANKING order="5" place="5" resultid="3576" />
                    <RANKING order="6" place="6" resultid="4808" />
                    <RANKING order="7" place="7" resultid="3404" />
                    <RANKING order="8" place="8" resultid="3338" />
                    <RANKING order="9" place="9" resultid="2252" />
                    <RANKING order="10" place="10" resultid="3917" />
                    <RANKING order="11" place="-1" resultid="3356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4317" />
                    <RANKING order="2" place="2" resultid="2482" />
                    <RANKING order="3" place="3" resultid="4393" />
                    <RANKING order="4" place="4" resultid="3558" />
                    <RANKING order="5" place="5" resultid="3457" />
                    <RANKING order="6" place="-1" resultid="3981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4202" />
                    <RANKING order="2" place="2" resultid="2776" />
                    <RANKING order="3" place="3" resultid="2050" />
                    <RANKING order="4" place="4" resultid="3827" />
                    <RANKING order="5" place="5" resultid="1763" />
                    <RANKING order="6" place="6" resultid="4325" />
                    <RANKING order="7" place="-1" resultid="2844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4332" />
                    <RANKING order="2" place="2" resultid="2681" />
                    <RANKING order="3" place="3" resultid="2427" />
                    <RANKING order="4" place="4" resultid="4657" />
                    <RANKING order="5" place="5" resultid="2284" />
                    <RANKING order="6" place="6" resultid="4339" />
                    <RANKING order="7" place="-1" resultid="2567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1235" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4032" />
                    <RANKING order="2" place="2" resultid="3727" />
                    <RANKING order="3" place="3" resultid="3807" />
                    <RANKING order="4" place="4" resultid="2246" />
                    <RANKING order="5" place="5" resultid="2093" />
                    <RANKING order="6" place="6" resultid="6033" />
                    <RANKING order="7" place="7" resultid="2899" />
                    <RANKING order="8" place="8" resultid="2834" />
                    <RANKING order="9" place="9" resultid="3041" />
                    <RANKING order="10" place="-1" resultid="2065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1236" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1857" />
                    <RANKING order="2" place="2" resultid="3769" />
                    <RANKING order="3" place="3" resultid="2105" />
                    <RANKING order="4" place="4" resultid="2830" />
                    <RANKING order="5" place="5" resultid="3222" />
                    <RANKING order="6" place="6" resultid="3963" />
                    <RANKING order="7" place="7" resultid="3002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3718" />
                    <RANKING order="2" place="2" resultid="4472" />
                    <RANKING order="3" place="3" resultid="3956" />
                    <RANKING order="4" place="4" resultid="3814" />
                    <RANKING order="5" place="5" resultid="3709" />
                    <RANKING order="6" place="6" resultid="4216" />
                    <RANKING order="7" place="7" resultid="4347" />
                    <RANKING order="8" place="8" resultid="3009" />
                    <RANKING order="9" place="9" resultid="6548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4185" />
                    <RANKING order="2" place="2" resultid="3942" />
                    <RANKING order="3" place="3" resultid="4367" />
                    <RANKING order="4" place="4" resultid="2199" />
                    <RANKING order="5" place="5" resultid="2813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4156" />
                    <RANKING order="2" place="2" resultid="3205" />
                    <RANKING order="3" place="3" resultid="3597" />
                    <RANKING order="4" place="4" resultid="3197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3697" />
                    <RANKING order="2" place="2" resultid="4721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6126" daytime="11:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6127" daytime="11:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6128" daytime="11:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6129" daytime="11:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6130" daytime="11:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6131" daytime="11:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6132" daytime="11:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6133" daytime="11:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6134" daytime="11:35" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6135" daytime="11:35" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6136" daytime="11:35" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6137" daytime="11:40" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6138" daytime="11:40" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6139" daytime="11:40" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1243" daytime="11:40" gender="F" number="12" order="15" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1244" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4485" />
                    <RANKING order="2" place="2" resultid="3663" />
                    <RANKING order="3" place="3" resultid="2338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2336" />
                    <RANKING order="2" place="2" resultid="4252" />
                    <RANKING order="3" place="-1" resultid="4732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1886" />
                    <RANKING order="2" place="2" resultid="2339" />
                    <RANKING order="3" place="-1" resultid="1723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4251" />
                    <RANKING order="2" place="2" resultid="3018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1249" agemax="-1" agemin="280" name="F: 280 lat i starsi" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6519" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6520" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1250" daytime="11:50" gender="M" number="13" order="17" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1251" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3073" />
                    <RANKING order="2" place="2" resultid="2669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4488" />
                    <RANKING order="2" place="2" resultid="4730" />
                    <RANKING order="3" place="3" resultid="2587" />
                    <RANKING order="4" place="4" resultid="3417" />
                    <RANKING order="5" place="5" resultid="3664" />
                    <RANKING order="6" place="6" resultid="3419" />
                    <RANKING order="7" place="7" resultid="3502" />
                    <RANKING order="8" place="8" resultid="3075" />
                    <RANKING order="9" place="9" resultid="3421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4118" />
                    <RANKING order="2" place="2" resultid="2328" />
                    <RANKING order="3" place="3" resultid="2588" />
                    <RANKING order="4" place="4" resultid="1807" />
                    <RANKING order="5" place="5" resultid="2330" />
                    <RANKING order="6" place="6" resultid="6026" />
                    <RANKING order="7" place="7" resultid="4487" />
                    <RANKING order="8" place="-1" resultid="4486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4735" />
                    <RANKING order="2" place="2" resultid="3740" />
                    <RANKING order="3" place="3" resultid="2589" />
                    <RANKING order="4" place="4" resultid="1891" />
                    <RANKING order="5" place="5" resultid="3020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1255" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4254" />
                    <RANKING order="2" place="2" resultid="3742" />
                    <RANKING order="3" place="3" resultid="3666" />
                    <RANKING order="4" place="4" resultid="3985" />
                    <RANKING order="5" place="5" resultid="4253" />
                    <RANKING order="6" place="6" resultid="2331" />
                    <RANKING order="7" place="7" resultid="6025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="-1" agemin="280" name="F: 280 lat i starsi" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1893" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6521" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6522" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6523" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6524" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6525" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6526" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1257" daytime="12:05" gender="F" number="14" order="19" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1258" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2647" />
                    <RANKING order="2" place="2" resultid="3924" />
                    <RANKING order="3" place="3" resultid="2027" />
                    <RANKING order="4" place="4" resultid="3626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3653" />
                    <RANKING order="2" place="2" resultid="3517" />
                    <RANKING order="3" place="3" resultid="2239" />
                    <RANKING order="4" place="4" resultid="4572" />
                    <RANKING order="5" place="5" resultid="4426" />
                    <RANKING order="6" place="6" resultid="1922" />
                    <RANKING order="7" place="7" resultid="4086" />
                    <RANKING order="8" place="8" resultid="4691" />
                    <RANKING order="9" place="9" resultid="4420" />
                    <RANKING order="10" place="10" resultid="2699" />
                    <RANKING order="11" place="-1" resultid="2278" />
                    <RANKING order="12" place="-1" resultid="2888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4684" />
                    <RANKING order="2" place="2" resultid="4598" />
                    <RANKING order="3" place="3" resultid="2036" />
                    <RANKING order="4" place="4" resultid="2827" />
                    <RANKING order="5" place="5" resultid="4056" />
                    <RANKING order="6" place="6" resultid="3513" />
                    <RANKING order="7" place="7" resultid="4448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3525" />
                    <RANKING order="2" place="2" resultid="4237" />
                    <RANKING order="3" place="3" resultid="4300" />
                    <RANKING order="4" place="4" resultid="4048" />
                    <RANKING order="5" place="5" resultid="4390" />
                    <RANKING order="6" place="6" resultid="3266" />
                    <RANKING order="7" place="7" resultid="2148" />
                    <RANKING order="8" place="8" resultid="3047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4196" />
                    <RANKING order="2" place="2" resultid="4413" />
                    <RANKING order="3" place="3" resultid="6549" />
                    <RANKING order="4" place="4" resultid="2881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2469" />
                    <RANKING order="2" place="2" resultid="2137" />
                    <RANKING order="3" place="3" resultid="4794" />
                    <RANKING order="4" place="4" resultid="4381" />
                    <RANKING order="5" place="5" resultid="2411" />
                    <RANKING order="6" place="6" resultid="4580" />
                    <RANKING order="7" place="7" resultid="2310" />
                    <RANKING order="8" place="8" resultid="4665" />
                    <RANKING order="9" place="-1" resultid="2560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1845" />
                    <RANKING order="2" place="2" resultid="2000" />
                    <RANKING order="3" place="3" resultid="1946" />
                    <RANKING order="4" place="4" resultid="1769" />
                    <RANKING order="5" place="5" resultid="3472" />
                    <RANKING order="6" place="6" resultid="3143" />
                    <RANKING order="7" place="-1" resultid="2738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2771" />
                    <RANKING order="2" place="2" resultid="3930" />
                    <RANKING order="3" place="3" resultid="1876" />
                    <RANKING order="4" place="4" resultid="4190" />
                    <RANKING order="5" place="5" resultid="2954" />
                    <RANKING order="6" place="6" resultid="4438" />
                    <RANKING order="7" place="7" resultid="2808" />
                    <RANKING order="8" place="8" resultid="2939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2946" />
                    <RANKING order="2" place="2" resultid="2932" />
                    <RANKING order="3" place="-1" resultid="4458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1269" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1270" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1271" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6148" daytime="12:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6149" daytime="12:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6150" daytime="12:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6151" daytime="12:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6152" daytime="12:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6153" daytime="12:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6154" daytime="12:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6155" daytime="12:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6156" daytime="12:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6157" daytime="12:25" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6158" daytime="12:25" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1272" daytime="12:30" gender="M" number="15" order="20" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1273" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2752" />
                    <RANKING order="2" place="2" resultid="2074" />
                    <RANKING order="3" place="3" resultid="3875" />
                    <RANKING order="4" place="4" resultid="2018" />
                    <RANKING order="5" place="5" resultid="4619" />
                    <RANKING order="6" place="6" resultid="2213" />
                    <RANKING order="7" place="7" resultid="3063" />
                    <RANKING order="8" place="8" resultid="2418" />
                    <RANKING order="9" place="9" resultid="4530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4633" />
                    <RANKING order="2" place="2" resultid="4539" />
                    <RANKING order="3" place="3" resultid="2082" />
                    <RANKING order="4" place="4" resultid="4313" />
                    <RANKING order="5" place="5" resultid="4433" />
                    <RANKING order="6" place="6" resultid="3860" />
                    <RANKING order="7" place="7" resultid="3786" />
                    <RANKING order="8" place="8" resultid="2583" />
                    <RANKING order="9" place="9" resultid="4105" />
                    <RANKING order="10" place="10" resultid="2115" />
                    <RANKING order="11" place="11" resultid="4093" />
                    <RANKING order="12" place="-1" resultid="4247" />
                    <RANKING order="13" place="-1" resultid="4698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3284" />
                    <RANKING order="2" place="2" resultid="3640" />
                    <RANKING order="3" place="3" resultid="4468" />
                    <RANKING order="4" place="4" resultid="4100" />
                    <RANKING order="5" place="5" resultid="3484" />
                    <RANKING order="6" place="6" resultid="3605" />
                    <RANKING order="7" place="7" resultid="1785" />
                    <RANKING order="8" place="8" resultid="3821" />
                    <RANKING order="9" place="9" resultid="4766" />
                    <RANKING order="10" place="10" resultid="3577" />
                    <RANKING order="11" place="11" resultid="3366" />
                    <RANKING order="12" place="12" resultid="3377" />
                    <RANKING order="13" place="13" resultid="3348" />
                    <RANKING order="14" place="14" resultid="4355" />
                    <RANKING order="15" place="15" resultid="3352" />
                    <RANKING order="16" place="16" resultid="2187" />
                    <RANKING order="17" place="17" resultid="4074" />
                    <RANKING order="18" place="18" resultid="3918" />
                    <RANKING order="19" place="-1" resultid="3291" />
                    <RANKING order="20" place="-1" resultid="3357" />
                    <RANKING order="21" place="-1" resultid="3373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2483" />
                    <RANKING order="2" place="2" resultid="3304" />
                    <RANKING order="3" place="3" resultid="4024" />
                    <RANKING order="4" place="4" resultid="4814" />
                    <RANKING order="5" place="5" resultid="2544" />
                    <RANKING order="6" place="6" resultid="2464" />
                    <RANKING order="7" place="7" resultid="3384" />
                    <RANKING order="8" place="8" resultid="3559" />
                    <RANKING order="9" place="9" resultid="2397" />
                    <RANKING order="10" place="10" resultid="2912" />
                    <RANKING order="11" place="11" resultid="4605" />
                    <RANKING order="12" place="12" resultid="1776" />
                    <RANKING order="13" place="-1" resultid="2438" />
                    <RANKING order="14" place="-1" resultid="2896" />
                    <RANKING order="15" place="-1" resultid="3489" />
                    <RANKING order="16" place="-1" resultid="4394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2823" />
                    <RANKING order="2" place="2" resultid="2777" />
                    <RANKING order="3" place="3" resultid="2190" />
                    <RANKING order="4" place="4" resultid="3168" />
                    <RANKING order="5" place="5" resultid="1751" />
                    <RANKING order="6" place="6" resultid="4203" />
                    <RANKING order="7" place="7" resultid="2522" />
                    <RANKING order="8" place="8" resultid="3892" />
                    <RANKING order="9" place="9" resultid="3230" />
                    <RANKING order="10" place="10" resultid="2043" />
                    <RANKING order="11" place="-1" resultid="2476" />
                    <RANKING order="12" place="-1" resultid="3244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3547" />
                    <RANKING order="2" place="2" resultid="3506" />
                    <RANKING order="3" place="3" resultid="2782" />
                    <RANKING order="4" place="4" resultid="1937" />
                    <RANKING order="5" place="5" resultid="2682" />
                    <RANKING order="6" place="6" resultid="4658" />
                    <RANKING order="7" place="7" resultid="3969" />
                    <RANKING order="8" place="8" resultid="2428" />
                    <RANKING order="9" place="9" resultid="4081" />
                    <RANKING order="10" place="10" resultid="3252" />
                    <RANKING order="11" place="11" resultid="3725" />
                    <RANKING order="12" place="12" resultid="2271" />
                    <RANKING order="13" place="13" resultid="4387" />
                    <RANKING order="14" place="-1" resultid="2169" />
                    <RANKING order="15" place="-1" resultid="2381" />
                    <RANKING order="16" place="-1" resultid="2694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4306" />
                    <RANKING order="2" place="2" resultid="2433" />
                    <RANKING order="3" place="3" resultid="2529" />
                    <RANKING order="4" place="4" resultid="4717" />
                    <RANKING order="5" place="5" resultid="3321" />
                    <RANKING order="6" place="6" resultid="4006" />
                    <RANKING order="7" place="7" resultid="2900" />
                    <RANKING order="8" place="8" resultid="1882" />
                    <RANKING order="9" place="9" resultid="2177" />
                    <RANKING order="10" place="10" resultid="4405" />
                    <RANKING order="11" place="-1" resultid="2066" />
                    <RANKING order="12" place="-1" resultid="2537" />
                    <RANKING order="13" place="-1" resultid="3496" />
                    <RANKING order="14" place="-1" resultid="4626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4361" />
                    <RANKING order="2" place="2" resultid="4142" />
                    <RANKING order="3" place="3" resultid="3735" />
                    <RANKING order="4" place="4" resultid="2058" />
                    <RANKING order="5" place="5" resultid="2760" />
                    <RANKING order="6" place="6" resultid="2106" />
                    <RANKING order="7" place="7" resultid="2765" />
                    <RANKING order="8" place="8" resultid="3055" />
                    <RANKING order="9" place="-1" resultid="3532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4473" />
                    <RANKING order="2" place="2" resultid="3719" />
                    <RANKING order="3" place="3" resultid="4671" />
                    <RANKING order="4" place="4" resultid="3584" />
                    <RANKING order="5" place="5" resultid="2982" />
                    <RANKING order="6" place="6" resultid="2122" />
                    <RANKING order="7" place="7" resultid="4348" />
                    <RANKING order="8" place="8" resultid="2619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2231" />
                    <RANKING order="2" place="2" resultid="2636" />
                    <RANKING order="3" place="3" resultid="1850" />
                    <RANKING order="4" place="4" resultid="4368" />
                    <RANKING order="5" place="-1" resultid="2974" />
                    <RANKING order="6" place="-1" resultid="3712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4157" />
                    <RANKING order="2" place="2" resultid="3598" />
                    <RANKING order="3" place="3" resultid="3198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3763" />
                    <RANKING order="2" place="2" resultid="1664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6515" agemax="89" agemin="85" name="M: 85 - 89 lat" />
                <AGEGROUP agegroupid="1286" agemax="-1" agemin="90" name="N: 90 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1864" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6159" daytime="12:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6160" daytime="12:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6161" daytime="12:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6162" daytime="12:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6163" daytime="12:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6164" daytime="12:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6165" daytime="12:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6166" daytime="12:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6167" daytime="12:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6168" daytime="12:50" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6169" daytime="12:50" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6170" daytime="12:50" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6171" daytime="12:55" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6172" daytime="12:55" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="6173" daytime="12:55" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="6174" daytime="12:55" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="6175" daytime="13:00" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="6176" daytime="13:00" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="6177" daytime="13:00" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="6178" daytime="13:05" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="6179" daytime="13:05" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="6180" daytime="13:05" number="22" order="22" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1287" daytime="13:10" gender="F" number="16" order="21" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1288" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1289" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="44" agemin="40" name="D: 40 - 44 lat" />
                <AGEGROUP agegroupid="1293" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3778" />
                    <RANKING order="2" place="2" resultid="1990" />
                    <RANKING order="3" place="3" resultid="1959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1297" agemax="69" agemin="65" name="I: 65 - 69 lat" />
                <AGEGROUP agegroupid="1298" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1299" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1300" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1301" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6181" daytime="13:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6182" daytime="13:15" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="13:20" gender="M" number="17" order="22" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1303" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4563" />
                    <RANKING order="2" place="2" resultid="2075" />
                    <RANKING order="3" place="3" resultid="2864" />
                    <RANKING order="4" place="4" resultid="4551" />
                    <RANKING order="5" place="-1" resultid="1734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4634" />
                    <RANKING order="2" place="2" resultid="2423" />
                    <RANKING order="3" place="3" resultid="2083" />
                    <RANKING order="4" place="4" resultid="3412" />
                    <RANKING order="5" place="-1" resultid="4094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4713" />
                    <RANKING order="2" place="2" resultid="3646" />
                    <RANKING order="3" place="3" resultid="2506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2491" />
                    <RANKING order="2" place="2" resultid="2257" />
                    <RANKING order="3" place="3" resultid="3180" />
                    <RANKING order="4" place="4" resultid="2499" />
                    <RANKING order="5" place="5" resultid="2552" />
                    <RANKING order="6" place="-1" resultid="2849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3128" />
                    <RANKING order="2" place="2" resultid="4232" />
                    <RANKING order="3" place="3" resultid="3121" />
                    <RANKING order="4" place="4" resultid="1743" />
                    <RANKING order="5" place="5" resultid="3828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3540" />
                    <RANKING order="2" place="2" resultid="2403" />
                    <RANKING order="3" place="3" resultid="2568" />
                    <RANKING order="4" place="4" resultid="1870" />
                    <RANKING order="5" place="-1" resultid="2675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4802" />
                    <RANKING order="2" place="2" resultid="2530" />
                    <RANKING order="3" place="3" resultid="1802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3705" />
                    <RANKING order="2" place="2" resultid="1858" />
                    <RANKING order="3" place="3" resultid="3846" />
                    <RANKING order="4" place="4" resultid="2714" />
                    <RANKING order="5" place="5" resultid="2918" />
                    <RANKING order="6" place="6" resultid="2907" />
                    <RANKING order="7" place="-1" resultid="1832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4672" />
                    <RANKING order="2" place="2" resultid="3214" />
                    <RANKING order="3" place="3" resultid="3911" />
                    <RANKING order="4" place="4" resultid="6541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2232" />
                    <RANKING order="2" place="2" resultid="1851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3206" />
                    <RANKING order="2" place="2" resultid="3158" />
                    <RANKING order="3" place="3" resultid="3854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1316" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6183" daytime="13:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6184" daytime="13:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6185" daytime="13:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6186" daytime="13:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6187" daytime="13:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6188" daytime="13:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6189" daytime="13:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6190" daytime="13:50" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6191" daytime="13:50" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2012-11-24" daytime="16:00" name="Blok III" number="3" warmupfrom="15:00">
          <EVENTS>
            <EVENT eventid="1318" daytime="16:00" gender="F" number="18" order="22" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1319" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2100" />
                    <RANKING order="2" place="2" resultid="2648" />
                    <RANKING order="3" place="3" resultid="2722" />
                    <RANKING order="4" place="4" resultid="3796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1320" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2279" />
                    <RANKING order="2" place="2" resultid="3312" />
                    <RANKING order="3" place="3" resultid="3654" />
                    <RANKING order="4" place="4" resultid="2209" />
                    <RANKING order="5" place="5" resultid="4573" />
                    <RANKING order="6" place="6" resultid="4692" />
                    <RANKING order="7" place="7" resultid="2461" />
                    <RANKING order="8" place="-1" resultid="2889" />
                    <RANKING order="9" place="-1" resultid="4087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1321" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4063" />
                    <RANKING order="2" place="2" resultid="2037" />
                    <RANKING order="3" place="3" resultid="4599" />
                    <RANKING order="4" place="4" resultid="3514" />
                    <RANKING order="5" place="-1" resultid="3634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1322" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3612" />
                    <RANKING order="2" place="2" resultid="3267" />
                    <RANKING order="3" place="3" resultid="3048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1323" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4480" />
                    <RANKING order="2" place="2" resultid="3260" />
                    <RANKING order="3" place="3" resultid="4113" />
                    <RANKING order="4" place="4" resultid="2882" />
                    <RANKING order="5" place="5" resultid="2262" />
                    <RANKING order="6" place="-1" resultid="4197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1324" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2132" />
                    <RANKING order="2" place="2" resultid="4382" />
                    <RANKING order="3" place="3" resultid="4581" />
                    <RANKING order="4" place="4" resultid="4453" />
                    <RANKING order="5" place="5" resultid="3521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1325" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1846" />
                    <RANKING order="2" place="2" resultid="2143" />
                    <RANKING order="3" place="3" resultid="2001" />
                    <RANKING order="4" place="4" resultid="4679" />
                    <RANKING order="5" place="5" resultid="1770" />
                    <RANKING order="6" place="6" resultid="3466" />
                    <RANKING order="7" place="7" resultid="3473" />
                    <RANKING order="8" place="8" resultid="2996" />
                    <RANKING order="9" place="9" resultid="3144" />
                    <RANKING order="10" place="-1" resultid="4229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1326" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3937" />
                    <RANKING order="2" place="2" resultid="3136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1327" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3931" />
                    <RANKING order="2" place="2" resultid="2156" />
                    <RANKING order="3" place="3" resultid="4138" />
                    <RANKING order="4" place="4" resultid="2940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1328" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4153" />
                    <RANKING order="2" place="2" resultid="4177" />
                    <RANKING order="3" place="3" resultid="4222" />
                    <RANKING order="4" place="4" resultid="2933" />
                    <RANKING order="5" place="5" resultid="2947" />
                    <RANKING order="6" place="6" resultid="2962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1329" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1815" />
                    <RANKING order="2" place="2" resultid="2969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1330" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6512" />
                    <RANKING order="2" place="2" resultid="4653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1331" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1332" agemax="-1" agemin="85" name="M: 85 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1979" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6192" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6193" daytime="16:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6194" daytime="16:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6195" daytime="16:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6196" daytime="16:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6197" daytime="16:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6198" daytime="16:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6199" daytime="16:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6200" daytime="16:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6201" daytime="16:15" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1333" daytime="16:15" gender="M" number="19" order="23" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1334" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2643" />
                    <RANKING order="2" place="2" resultid="4535" />
                    <RANKING order="3" place="2" resultid="4564" />
                    <RANKING order="4" place="4" resultid="3064" />
                    <RANKING order="5" place="5" resultid="3794" />
                    <RANKING order="6" place="-1" resultid="1735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1335" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4556" />
                    <RANKING order="2" place="2" resultid="4464" />
                    <RANKING order="3" place="3" resultid="2726" />
                    <RANKING order="4" place="4" resultid="3398" />
                    <RANKING order="5" place="5" resultid="2652" />
                    <RANKING order="6" place="6" resultid="2116" />
                    <RANKING order="7" place="7" resultid="2584" />
                    <RANKING order="8" place="8" resultid="3392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1336" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4709" />
                    <RANKING order="2" place="2" resultid="3362" />
                    <RANKING order="3" place="3" resultid="1790" />
                    <RANKING order="4" place="4" resultid="4809" />
                    <RANKING order="5" place="5" resultid="3578" />
                    <RANKING order="6" place="6" resultid="3339" />
                    <RANKING order="7" place="7" resultid="3345" />
                    <RANKING order="8" place="8" resultid="2459" />
                    <RANKING order="9" place="9" resultid="3919" />
                    <RANKING order="10" place="-1" resultid="3097" />
                    <RANKING order="11" place="-1" resultid="3236" />
                    <RANKING order="12" place="-1" resultid="3374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1337" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2577" />
                    <RANKING order="2" place="2" resultid="2545" />
                    <RANKING order="3" place="3" resultid="2500" />
                    <RANKING order="4" place="4" resultid="2316" />
                    <RANKING order="5" place="-1" resultid="3492" />
                    <RANKING order="6" place="-1" resultid="4025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1338" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3869" />
                    <RANKING order="2" place="2" resultid="3450" />
                    <RANKING order="3" place="3" resultid="2226" />
                    <RANKING order="4" place="4" resultid="2729" />
                    <RANKING order="5" place="5" resultid="3975" />
                    <RANKING order="6" place="6" resultid="2442" />
                    <RANKING order="7" place="7" resultid="4326" />
                    <RANKING order="8" place="-1" resultid="2845" />
                    <RANKING order="9" place="-1" resultid="3245" />
                    <RANKING order="10" place="-1" resultid="4012" />
                    <RANKING order="11" place="-1" resultid="4015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1339" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3507" />
                    <RANKING order="2" place="2" resultid="2783" />
                    <RANKING order="3" place="3" resultid="3970" />
                    <RANKING order="4" place="4" resultid="2170" />
                    <RANKING order="5" place="5" resultid="4340" />
                    <RANKING order="6" place="6" resultid="3715" />
                    <RANKING order="7" place="-1" resultid="3884" />
                    <RANKING order="8" place="-1" resultid="2382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1340" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4627" />
                    <RANKING order="2" place="2" resultid="3553" />
                    <RANKING order="3" place="3" resultid="2538" />
                    <RANKING order="4" place="4" resultid="4776" />
                    <RANKING order="5" place="5" resultid="1883" />
                    <RANKING order="6" place="6" resultid="4774" />
                    <RANKING order="7" place="7" resultid="2178" />
                    <RANKING order="8" place="8" resultid="4406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1341" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2745" />
                    <RANKING order="2" place="2" resultid="1795" />
                    <RANKING order="3" place="3" resultid="2831" />
                    <RANKING order="4" place="4" resultid="2766" />
                    <RANKING order="5" place="5" resultid="3660" />
                    <RANKING order="6" place="6" resultid="1833" />
                    <RANKING order="7" place="7" resultid="3731" />
                    <RANKING order="8" place="8" resultid="3003" />
                    <RANKING order="9" place="9" resultid="2919" />
                    <RANKING order="10" place="10" resultid="3056" />
                    <RANKING order="11" place="11" resultid="3152" />
                    <RANKING order="12" place="12" resultid="2908" />
                    <RANKING order="13" place="13" resultid="2289" />
                    <RANKING order="14" place="-1" resultid="4068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1342" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4589" />
                    <RANKING order="2" place="2" resultid="3774" />
                    <RANKING order="3" place="3" resultid="1828" />
                    <RANKING order="4" place="4" resultid="1953" />
                    <RANKING order="5" place="5" resultid="3571" />
                    <RANKING order="6" place="6" resultid="4241" />
                    <RANKING order="7" place="7" resultid="2302" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1343" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3950" />
                    <RANKING order="2" place="2" resultid="2689" />
                    <RANKING order="3" place="3" resultid="4369" />
                    <RANKING order="4" place="4" resultid="2989" />
                    <RANKING order="5" place="5" resultid="2814" />
                    <RANKING order="6" place="-1" resultid="2975" />
                    <RANKING order="7" place="-1" resultid="3713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4158" />
                    <RANKING order="2" place="2" resultid="4182" />
                    <RANKING order="3" place="3" resultid="3159" />
                    <RANKING order="4" place="4" resultid="1983" />
                    <RANKING order="5" place="5" resultid="3199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3699" />
                    <RANKING order="2" place="2" resultid="4293" />
                    <RANKING order="3" place="-1" resultid="4722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1347" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6202" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6203" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6204" daytime="16:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6205" daytime="16:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6206" daytime="16:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6207" daytime="16:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6208" daytime="16:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6209" daytime="16:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6210" daytime="16:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6211" daytime="16:30" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6212" daytime="16:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6213" daytime="16:30" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6214" daytime="16:30" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6215" daytime="16:30" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="6216" daytime="16:35" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="6217" daytime="16:35" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1348" daytime="16:35" gender="F" number="20" order="24" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1349" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2305" />
                    <RANKING order="2" place="2" resultid="4737" />
                    <RANKING order="3" place="3" resultid="2706" />
                    <RANKING order="4" place="4" resultid="2449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1350" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3313" />
                    <RANKING order="2" place="2" resultid="3518" />
                    <RANKING order="3" place="3" resultid="4427" />
                    <RANKING order="4" place="4" resultid="4088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1351" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2857" />
                    <RANKING order="2" place="2" resultid="2390" />
                    <RANKING order="3" place="3" resultid="3479" />
                    <RANKING order="4" place="4" resultid="2194" />
                    <RANKING order="5" place="-1" resultid="4685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4238" />
                    <RANKING order="2" place="2" resultid="3526" />
                    <RANKING order="3" place="3" resultid="2149" />
                    <RANKING order="4" place="-1" resultid="2840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1353" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3802" />
                    <RANKING order="2" place="2" resultid="2138" />
                    <RANKING order="3" place="3" resultid="2561" />
                    <RANKING order="4" place="4" resultid="4666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1355" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1840" />
                    <RANKING order="2" place="2" resultid="3779" />
                    <RANKING order="3" place="3" resultid="2002" />
                    <RANKING order="4" place="4" resultid="3619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1356" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2221" />
                    <RANKING order="2" place="2" resultid="1823" />
                    <RANKING order="3" place="3" resultid="1974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1357" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4167" />
                    <RANKING order="2" place="2" resultid="1877" />
                    <RANKING order="3" place="3" resultid="2955" />
                    <RANKING order="4" place="4" resultid="1967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1358" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4173" />
                    <RANKING order="2" place="2" resultid="2162" />
                    <RANKING order="3" place="3" resultid="2963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1359" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1360" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1361" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1362" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6218" daytime="16:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6219" daytime="16:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6220" daytime="16:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6221" daytime="16:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6222" daytime="16:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6223" daytime="16:45" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1363" daytime="16:45" gender="M" number="21" order="25" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1364" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2801" />
                    <RANKING order="2" place="2" resultid="2019" />
                    <RANKING order="3" place="3" resultid="2076" />
                    <RANKING order="4" place="4" resultid="4620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1365" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3101" />
                    <RANKING order="2" place="2" resultid="4635" />
                    <RANKING order="3" place="3" resultid="4699" />
                    <RANKING order="4" place="4" resultid="4314" />
                    <RANKING order="5" place="5" resultid="3861" />
                    <RANKING order="6" place="6" resultid="4434" />
                    <RANKING order="7" place="7" resultid="2084" />
                    <RANKING order="8" place="8" resultid="3413" />
                    <RANKING order="9" place="9" resultid="4465" />
                    <RANKING order="10" place="10" resultid="3787" />
                    <RANKING order="11" place="11" resultid="4095" />
                    <RANKING order="12" place="12" resultid="4106" />
                    <RANKING order="13" place="-1" resultid="3461" />
                    <RANKING order="14" place="-1" resultid="3071" />
                    <RANKING order="15" place="-1" resultid="4248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1366" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4444" />
                    <RANKING order="2" place="2" resultid="4710" />
                    <RANKING order="3" place="3" resultid="3485" />
                    <RANKING order="4" place="4" resultid="1786" />
                    <RANKING order="5" place="5" resultid="4101" />
                    <RANKING order="6" place="6" resultid="4714" />
                    <RANKING order="7" place="7" resultid="3367" />
                    <RANKING order="8" place="8" resultid="3363" />
                    <RANKING order="9" place="9" resultid="4075" />
                    <RANKING order="10" place="10" resultid="3353" />
                    <RANKING order="11" place="11" resultid="3349" />
                    <RANKING order="12" place="12" resultid="3378" />
                    <RANKING order="13" place="13" resultid="3647" />
                    <RANKING order="14" place="14" resultid="3565" />
                    <RANKING order="15" place="15" resultid="3405" />
                    <RANKING order="16" place="16" resultid="3237" />
                    <RANKING order="17" place="17" resultid="2507" />
                    <RANKING order="18" place="-1" resultid="3094" />
                    <RANKING order="19" place="-1" resultid="4245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1367" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4318" />
                    <RANKING order="2" place="2" resultid="4026" />
                    <RANKING order="3" place="3" resultid="4815" />
                    <RANKING order="4" place="4" resultid="3385" />
                    <RANKING order="5" place="5" resultid="3560" />
                    <RANKING order="6" place="6" resultid="2850" />
                    <RANKING order="7" place="7" resultid="4395" />
                    <RANKING order="8" place="8" resultid="2258" />
                    <RANKING order="9" place="9" resultid="2484" />
                    <RANKING order="10" place="10" resultid="4606" />
                    <RANKING order="11" place="-1" resultid="3982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1368" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2824" />
                    <RANKING order="2" place="2" resultid="2778" />
                    <RANKING order="3" place="3" resultid="3129" />
                    <RANKING order="4" place="4" resultid="2227" />
                    <RANKING order="5" place="5" resultid="2191" />
                    <RANKING order="6" place="6" resultid="3870" />
                    <RANKING order="7" place="7" resultid="2183" />
                    <RANKING order="8" place="8" resultid="4233" />
                    <RANKING order="9" place="9" resultid="1752" />
                    <RANKING order="10" place="10" resultid="1997" />
                    <RANKING order="11" place="11" resultid="3122" />
                    <RANKING order="12" place="12" resultid="3231" />
                    <RANKING order="13" place="13" resultid="1744" />
                    <RANKING order="14" place="14" resultid="3893" />
                    <RANKING order="15" place="15" resultid="3976" />
                    <RANKING order="16" place="-1" resultid="2443" />
                    <RANKING order="17" place="-1" resultid="4016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1369" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3508" />
                    <RANKING order="2" place="2" resultid="2683" />
                    <RANKING order="3" place="3" resultid="1938" />
                    <RANKING order="4" place="4" resultid="2569" />
                    <RANKING order="5" place="5" resultid="4082" />
                    <RANKING order="6" place="6" resultid="3253" />
                    <RANKING order="7" place="7" resultid="2404" />
                    <RANKING order="8" place="8" resultid="2285" />
                    <RANKING order="9" place="-1" resultid="2272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1370" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4307" />
                    <RANKING order="2" place="2" resultid="3808" />
                    <RANKING order="3" place="3" resultid="2247" />
                    <RANKING order="4" place="4" resultid="4718" />
                    <RANKING order="5" place="5" resultid="1803" />
                    <RANKING order="6" place="6" resultid="2901" />
                    <RANKING order="7" place="-1" resultid="3886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1371" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1796" />
                    <RANKING order="2" place="2" resultid="1859" />
                    <RANKING order="3" place="3" resultid="2746" />
                    <RANKING order="4" place="4" resultid="3706" />
                    <RANKING order="5" place="5" resultid="3736" />
                    <RANKING order="6" place="6" resultid="2059" />
                    <RANKING order="7" place="7" resultid="3847" />
                    <RANKING order="8" place="8" resultid="3004" />
                    <RANKING order="9" place="9" resultid="2909" />
                    <RANKING order="10" place="-1" resultid="4069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1372" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3585" />
                    <RANKING order="2" place="2" resultid="4349" />
                    <RANKING order="3" place="3" resultid="4217" />
                    <RANKING order="4" place="4" resultid="3815" />
                    <RANKING order="5" place="5" resultid="2620" />
                    <RANKING order="6" place="6" resultid="3010" />
                    <RANKING order="7" place="-1" resultid="4673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1373" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2637" />
                    <RANKING order="2" place="2" resultid="1852" />
                    <RANKING order="3" place="3" resultid="2205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1374" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3160" />
                    <RANKING order="2" place="2" resultid="3855" />
                    <RANKING order="3" place="3" resultid="3207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1375" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1376" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1377" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6224" daytime="16:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6225" daytime="16:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6226" daytime="16:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6227" daytime="16:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6228" daytime="16:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6229" daytime="16:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6230" daytime="16:50" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6231" daytime="16:55" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6232" daytime="16:55" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6233" daytime="16:55" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6234" daytime="16:55" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6235" daytime="16:55" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6236" daytime="17:00" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6237" daytime="17:00" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="6238" daytime="17:00" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="6239" daytime="17:00" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="6240" daytime="17:00" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="6241" daytime="17:05" number="18" order="18" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1378" daytime="17:05" gender="F" number="22" order="26" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1379" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2707" />
                    <RANKING order="2" place="2" resultid="2028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1380" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2240" />
                    <RANKING order="2" place="2" resultid="4041" />
                    <RANKING order="3" place="3" resultid="4693" />
                    <RANKING order="4" place="-1" resultid="3314" />
                    <RANKING order="5" place="-1" resultid="1923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1381" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3635" />
                    <RANKING order="2" place="2" resultid="2391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1382" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4301" />
                    <RANKING order="2" place="2" resultid="3997" />
                    <RANKING order="3" place="3" resultid="4049" />
                    <RANKING order="4" place="-1" resultid="4391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1383" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4210" />
                    <RANKING order="2" place="2" resultid="2294" />
                    <RANKING order="3" place="3" resultid="4114" />
                    <RANKING order="4" place="4" resultid="3297" />
                    <RANKING order="5" place="5" resultid="2263" />
                    <RANKING order="6" place="6" resultid="2883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1384" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2133" />
                    <RANKING order="2" place="2" resultid="2412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1385" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3838" />
                    <RANKING order="2" place="2" resultid="1991" />
                    <RANKING order="3" place="3" resultid="1771" />
                    <RANKING order="4" place="4" resultid="3620" />
                    <RANKING order="5" place="5" resultid="2997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1386" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3938" />
                    <RANKING order="2" place="2" resultid="4148" />
                    <RANKING order="3" place="3" resultid="3137" />
                    <RANKING order="4" place="4" resultid="2925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1387" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2772" />
                    <RANKING order="2" place="2" resultid="2941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1388" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1389" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4642" />
                    <RANKING order="2" place="-1" resultid="1816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1390" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4400" />
                    <RANKING order="2" place="2" resultid="4654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1391" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1392" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6242" daytime="17:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6243" daytime="17:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6244" daytime="17:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6245" daytime="17:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6246" daytime="17:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6247" daytime="17:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6248" daytime="17:20" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1393" daytime="17:25" gender="M" number="23" order="27" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1394" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2753" />
                    <RANKING order="2" place="2" resultid="2865" />
                    <RANKING order="3" place="3" resultid="4614" />
                    <RANKING order="4" place="4" resultid="4546" />
                    <RANKING order="5" place="5" resultid="4531" />
                    <RANKING order="6" place="-1" resultid="2656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1395" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3110" />
                    <RANKING order="2" place="2" resultid="2630" />
                    <RANKING order="3" place="3" resultid="3393" />
                    <RANKING order="4" place="-1" resultid="2735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1396" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3285" />
                    <RANKING order="2" place="2" resultid="3641" />
                    <RANKING order="3" place="3" resultid="3606" />
                    <RANKING order="4" place="4" resultid="2090" />
                    <RANKING order="5" place="5" resultid="3331" />
                    <RANKING order="6" place="6" resultid="3340" />
                    <RANKING order="7" place="7" resultid="3406" />
                    <RANKING order="8" place="8" resultid="3566" />
                    <RANKING order="9" place="9" resultid="2253" />
                    <RANKING order="10" place="10" resultid="3920" />
                    <RANKING order="11" place="-1" resultid="3358" />
                    <RANKING order="12" place="-1" resultid="3579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4319" />
                    <RANKING order="2" place="2" resultid="2485" />
                    <RANKING order="3" place="3" resultid="4396" />
                    <RANKING order="4" place="4" resultid="3561" />
                    <RANKING order="5" place="5" resultid="2553" />
                    <RANKING order="6" place="6" resultid="3458" />
                    <RANKING order="7" place="7" resultid="2873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1398" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4204" />
                    <RANKING order="2" place="2" resultid="2051" />
                    <RANKING order="3" place="3" resultid="3015" />
                    <RANKING order="4" place="4" resultid="2523" />
                    <RANKING order="5" place="5" resultid="3829" />
                    <RANKING order="6" place="6" resultid="1764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1399" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4333" />
                    <RANKING order="2" place="2" resultid="4659" />
                    <RANKING order="3" place="3" resultid="2429" />
                    <RANKING order="4" place="4" resultid="2570" />
                    <RANKING order="5" place="5" resultid="4772" />
                    <RANKING order="6" place="6" resultid="4341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1400" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4033" />
                    <RANKING order="2" place="2" resultid="3728" />
                    <RANKING order="3" place="3" resultid="3809" />
                    <RANKING order="4" place="4" resultid="2094" />
                    <RANKING order="5" place="5" resultid="6034" />
                    <RANKING order="6" place="6" resultid="3042" />
                    <RANKING order="7" place="7" resultid="4407" />
                    <RANKING order="8" place="-1" resultid="2248" />
                    <RANKING order="9" place="-1" resultid="2067" />
                    <RANKING order="10" place="-1" resultid="4770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1401" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4362" />
                    <RANKING order="2" place="2" resultid="3770" />
                    <RANKING order="3" place="3" resultid="3533" />
                    <RANKING order="4" place="4" resultid="2715" />
                    <RANKING order="5" place="5" resultid="3964" />
                    <RANKING order="6" place="6" resultid="2107" />
                    <RANKING order="7" place="7" resultid="3223" />
                    <RANKING order="8" place="8" resultid="3737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1402" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4474" />
                    <RANKING order="2" place="2" resultid="3720" />
                    <RANKING order="3" place="3" resultid="2515" />
                    <RANKING order="4" place="4" resultid="3957" />
                    <RANKING order="5" place="5" resultid="3912" />
                    <RANKING order="6" place="6" resultid="3710" />
                    <RANKING order="7" place="7" resultid="3572" />
                    <RANKING order="8" place="8" resultid="6542" />
                    <RANKING order="9" place="9" resultid="3011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1403" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4186" />
                    <RANKING order="2" place="2" resultid="3943" />
                    <RANKING order="3" place="3" resultid="3951" />
                    <RANKING order="4" place="4" resultid="2815" />
                    <RANKING order="5" place="-1" resultid="2200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1404" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3599" />
                    <RANKING order="2" place="2" resultid="6546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1405" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3700" />
                    <RANKING order="2" place="2" resultid="4723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1406" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                    <RANKING order="2" place="2" resultid="3693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1407" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6249" daytime="17:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6250" daytime="17:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6251" daytime="17:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6252" daytime="17:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6253" daytime="17:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6254" daytime="17:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6255" daytime="17:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6256" daytime="17:40" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6257" daytime="17:40" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6258" daytime="17:45" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6259" daytime="17:45" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6260" daytime="17:45" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6261" daytime="17:50" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6262" daytime="17:50" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1408" daytime="17:50" gender="F" number="24" order="29" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1409" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1410" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4489" />
                    <RANKING order="2" place="2" resultid="3662" />
                    <RANKING order="3" place="3" resultid="2337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1411" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4256" />
                    <RANKING order="2" place="2" resultid="2335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1412" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2334" />
                    <RANKING order="2" place="2" resultid="1888" />
                    <RANKING order="3" place="3" resultid="1724" />
                    <RANKING order="4" place="4" resultid="4731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1413" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4255" />
                    <RANKING order="2" place="2" resultid="3019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1414" agemax="-1" agemin="280" name="F: 280 lat i starsi" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6527" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6528" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1415" daytime="18:00" gender="M" number="25" order="30" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1416" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1417" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4729" />
                    <RANKING order="2" place="2" resultid="4490" />
                    <RANKING order="3" place="3" resultid="3665" />
                    <RANKING order="4" place="4" resultid="3418" />
                    <RANKING order="5" place="5" resultid="2590" />
                    <RANKING order="6" place="6" resultid="3420" />
                    <RANKING order="7" place="7" resultid="3422" />
                    <RANKING order="8" place="8" resultid="6518" />
                    <RANKING order="9" place="9" resultid="3076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1418" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4120" />
                    <RANKING order="2" place="2" resultid="2332" />
                    <RANKING order="3" place="3" resultid="2591" />
                    <RANKING order="4" place="4" resultid="4491" />
                    <RANKING order="5" place="5" resultid="2329" />
                    <RANKING order="6" place="6" resultid="6027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4736" />
                    <RANKING order="2" place="2" resultid="3741" />
                    <RANKING order="3" place="3" resultid="4777" />
                    <RANKING order="4" place="4" resultid="2592" />
                    <RANKING order="5" place="5" resultid="1892" />
                    <RANKING order="6" place="6" resultid="4258" />
                    <RANKING order="7" place="7" resultid="4492" />
                    <RANKING order="8" place="-1" resultid="3021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1420" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4257" />
                    <RANKING order="2" place="2" resultid="3743" />
                    <RANKING order="3" place="3" resultid="3667" />
                    <RANKING order="4" place="4" resultid="2333" />
                    <RANKING order="5" place="-1" resultid="3271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1421" agemax="-1" agemin="280" name="F: 280 lat i starsi" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1894" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6529" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6530" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6531" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6532" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6533" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6534" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1422" daytime="18:10" gender="F" number="26" order="31" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1423" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3925" />
                    <RANKING order="2" place="2" resultid="2029" />
                    <RANKING order="3" place="-1" resultid="3627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1424" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4574" />
                    <RANKING order="2" place="2" resultid="1924" />
                    <RANKING order="3" place="3" resultid="4421" />
                    <RANKING order="4" place="4" resultid="2700" />
                    <RANKING order="5" place="-1" resultid="2890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2858" />
                    <RANKING order="2" place="2" resultid="4600" />
                    <RANKING order="3" place="3" resultid="4057" />
                    <RANKING order="4" place="4" resultid="3480" />
                    <RANKING order="5" place="5" resultid="2195" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1658" />
                    <RANKING order="2" place="2" resultid="3527" />
                    <RANKING order="3" place="3" resultid="4050" />
                    <RANKING order="4" place="4" resultid="2150" />
                    <RANKING order="5" place="5" resultid="3049" />
                    <RANKING order="6" place="-1" resultid="3268" />
                    <RANKING order="7" place="-1" resultid="4302" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4414" />
                    <RANKING order="2" place="2" resultid="3261" />
                    <RANKING order="3" place="3" resultid="3298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1428" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2470" />
                    <RANKING order="2" place="2" resultid="4795" />
                    <RANKING order="3" place="3" resultid="4383" />
                    <RANKING order="4" place="4" resultid="2413" />
                    <RANKING order="5" place="5" resultid="2311" />
                    <RANKING order="6" place="6" resultid="4454" />
                    <RANKING order="7" place="7" resultid="4667" />
                    <RANKING order="8" place="-1" resultid="4582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1429" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1947" />
                    <RANKING order="2" place="2" resultid="3145" />
                    <RANKING order="3" place="-1" resultid="2739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1824" />
                    <RANKING order="2" place="2" resultid="1975" />
                    <RANKING order="3" place="3" resultid="2926" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1431" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4191" />
                    <RANKING order="2" place="2" resultid="2956" />
                    <RANKING order="3" place="3" resultid="4439" />
                    <RANKING order="4" place="4" resultid="2809" />
                    <RANKING order="5" place="-1" resultid="3932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1432" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2163" />
                    <RANKING order="2" place="2" resultid="2934" />
                    <RANKING order="3" place="-1" resultid="4459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1433" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1434" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1435" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1436" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6270" daytime="18:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6271" daytime="18:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6272" daytime="18:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6273" daytime="18:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6274" daytime="18:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6275" daytime="18:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6276" daytime="18:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6277" daytime="18:50" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1437" daytime="18:50" gender="M" number="27" order="32" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1438" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3876" />
                    <RANKING order="2" place="2" resultid="2077" />
                    <RANKING order="3" place="3" resultid="2214" />
                    <RANKING order="4" place="4" resultid="4621" />
                    <RANKING order="5" place="5" resultid="3888" />
                    <RANKING order="6" place="-1" resultid="2802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1439" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4636" />
                    <RANKING order="2" place="2" resultid="2085" />
                    <RANKING order="3" place="3" resultid="3904" />
                    <RANKING order="4" place="4" resultid="2424" />
                    <RANKING order="5" place="5" resultid="3788" />
                    <RANKING order="6" place="6" resultid="4107" />
                    <RANKING order="7" place="7" resultid="4096" />
                    <RANKING order="8" place="8" resultid="2585" />
                    <RANKING order="9" place="-1" resultid="4540" />
                    <RANKING order="10" place="-1" resultid="4700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1440" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3286" />
                    <RANKING order="2" place="2" resultid="3642" />
                    <RANKING order="3" place="3" resultid="3822" />
                    <RANKING order="4" place="4" resultid="1782" />
                    <RANKING order="5" place="5" resultid="3379" />
                    <RANKING order="6" place="6" resultid="3368" />
                    <RANKING order="7" place="7" resultid="4356" />
                    <RANKING order="8" place="-1" resultid="3607" />
                    <RANKING order="9" place="-1" resultid="3648" />
                    <RANKING order="10" place="-1" resultid="4076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1441" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2492" />
                    <RANKING order="2" place="2" resultid="3305" />
                    <RANKING order="3" place="3" resultid="2546" />
                    <RANKING order="4" place="4" resultid="2465" />
                    <RANKING order="5" place="5" resultid="3386" />
                    <RANKING order="6" place="6" resultid="3115" />
                    <RANKING order="7" place="7" resultid="2913" />
                    <RANKING order="8" place="8" resultid="1777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3169" />
                    <RANKING order="2" place="2" resultid="4205" />
                    <RANKING order="3" place="3" resultid="1753" />
                    <RANKING order="4" place="4" resultid="2779" />
                    <RANKING order="5" place="5" resultid="2477" />
                    <RANKING order="6" place="6" resultid="2044" />
                    <RANKING order="7" place="7" resultid="4327" />
                    <RANKING order="8" place="-1" resultid="3246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4375" />
                    <RANKING order="2" place="2" resultid="3548" />
                    <RANKING order="3" place="3" resultid="2784" />
                    <RANKING order="4" place="4" resultid="4660" />
                    <RANKING order="5" place="5" resultid="2405" />
                    <RANKING order="6" place="6" resultid="2273" />
                    <RANKING order="7" place="-1" resultid="2383" />
                    <RANKING order="8" place="-1" resultid="2676" />
                    <RANKING order="9" place="-1" resultid="2695" />
                    <RANKING order="10" place="-1" resultid="3971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4803" />
                    <RANKING order="2" place="2" resultid="2434" />
                    <RANKING order="3" place="3" resultid="4007" />
                    <RANKING order="4" place="4" resultid="2179" />
                    <RANKING order="5" place="-1" resultid="2531" />
                    <RANKING order="6" place="-1" resultid="2902" />
                    <RANKING order="7" place="-1" resultid="2068" />
                    <RANKING order="8" place="-1" resultid="3322" />
                    <RANKING order="9" place="-1" resultid="4308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2761" />
                    <RANKING order="2" place="2" resultid="3848" />
                    <RANKING order="3" place="3" resultid="4143" />
                    <RANKING order="4" place="4" resultid="3707" />
                    <RANKING order="5" place="5" resultid="2060" />
                    <RANKING order="6" place="6" resultid="3534" />
                    <RANKING order="7" place="7" resultid="3057" />
                    <RANKING order="8" place="-1" resultid="3224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1446" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4475" />
                    <RANKING order="2" place="2" resultid="3721" />
                    <RANKING order="3" place="3" resultid="4674" />
                    <RANKING order="4" place="4" resultid="2123" />
                    <RANKING order="5" place="5" resultid="2983" />
                    <RANKING order="6" place="6" resultid="3215" />
                    <RANKING order="7" place="7" resultid="6543" />
                    <RANKING order="8" place="8" resultid="4350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2233" />
                    <RANKING order="2" place="2" resultid="4370" />
                    <RANKING order="3" place="3" resultid="2990" />
                    <RANKING order="4" place="-1" resultid="2201" />
                    <RANKING order="5" place="-1" resultid="2976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1448" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4159" />
                    <RANKING order="2" place="2" resultid="3600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1449" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3765" />
                    <RANKING order="2" place="2" resultid="1666" />
                    <RANKING order="3" place="3" resultid="2625" />
                    <RANKING order="4" place="4" resultid="3694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6516" agemax="89" agemin="85" name="M: 85 lat i starsi" />
                <AGEGROUP agegroupid="1451" agemax="-1" agemin="90" name="N: 90 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1865" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6278" daytime="18:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6279" daytime="19:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6280" daytime="19:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6281" daytime="19:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6282" daytime="19:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6283" daytime="19:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6284" daytime="19:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6285" daytime="19:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6286" daytime="19:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6287" daytime="19:25" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6288" daytime="19:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6289" daytime="19:30" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6290" daytime="19:35" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6291" daytime="19:35" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="6292" daytime="19:40" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1452" daytime="19:45" gender="F" number="28" order="33" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1453" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2101" />
                    <RANKING order="2" place="2" resultid="2450" />
                    <RANKING order="3" place="3" resultid="3628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1454" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3655" />
                    <RANKING order="2" place="2" resultid="4042" />
                    <RANKING order="3" place="3" resultid="2241" />
                    <RANKING order="4" place="4" resultid="4428" />
                    <RANKING order="5" place="5" resultid="4422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1455" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2038" />
                    <RANKING order="2" place="2" resultid="4058" />
                    <RANKING order="3" place="3" resultid="4449" />
                    <RANKING order="4" place="-1" resultid="4686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1456" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3613" />
                    <RANKING order="2" place="2" resultid="2793" />
                    <RANKING order="3" place="3" resultid="3998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1457" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4198" />
                    <RANKING order="2" place="2" resultid="4211" />
                    <RANKING order="3" place="3" resultid="2295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1458" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2139" />
                    <RANKING order="2" place="2" resultid="2562" />
                    <RANKING order="3" place="3" resultid="4796" />
                    <RANKING order="4" place="-1" resultid="3803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3839" />
                    <RANKING order="2" place="2" resultid="3780" />
                    <RANKING order="3" place="3" resultid="3474" />
                    <RANKING order="4" place="4" resultid="4680" />
                    <RANKING order="5" place="5" resultid="3467" />
                    <RANKING order="6" place="-1" resultid="1960" />
                    <RANKING order="7" place="-1" resultid="1992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1460" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1461" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4168" />
                    <RANKING order="2" place="2" resultid="2157" />
                    <RANKING order="3" place="3" resultid="1968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1462" agemax="69" agemin="65" name="I: 65 - 69 lat" />
                <AGEGROUP agegroupid="1463" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1464" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1465" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1466" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6293" daytime="19:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6294" daytime="19:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6295" daytime="19:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6296" daytime="19:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6297" daytime="20:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6298" daytime="20:05" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1467" daytime="20:05" gender="M" number="29" order="34" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1468" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2754" />
                    <RANKING order="2" place="2" resultid="4565" />
                    <RANKING order="3" place="3" resultid="2020" />
                    <RANKING order="4" place="4" resultid="4615" />
                    <RANKING order="5" place="5" resultid="3065" />
                    <RANKING order="6" place="-1" resultid="1736" />
                    <RANKING order="7" place="-1" resultid="2866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1469" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2659" />
                    <RANKING order="2" place="2" resultid="3399" />
                    <RANKING order="3" place="3" resultid="2663" />
                    <RANKING order="4" place="-1" resultid="3414" />
                    <RANKING order="5" place="-1" resultid="4557" />
                    <RANKING order="6" place="-1" resultid="3905" />
                    <RANKING order="7" place="-1" resultid="2667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1470" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3332" />
                    <RANKING order="2" place="2" resultid="2508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1471" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2493" />
                    <RANKING order="2" place="2" resultid="2578" />
                    <RANKING order="3" place="3" resultid="4816" />
                    <RANKING order="4" place="4" resultid="3181" />
                    <RANKING order="5" place="5" resultid="2554" />
                    <RANKING order="6" place="6" resultid="4607" />
                    <RANKING order="7" place="7" resultid="2869" />
                    <RANKING order="8" place="-1" resultid="2501" />
                    <RANKING order="9" place="-1" resultid="2851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1472" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3451" />
                    <RANKING order="2" place="2" resultid="2052" />
                    <RANKING order="3" place="3" resultid="2478" />
                    <RANKING order="4" place="4" resultid="2524" />
                    <RANKING order="5" place="5" resultid="3830" />
                    <RANKING order="6" place="6" resultid="3123" />
                    <RANKING order="7" place="7" resultid="1745" />
                    <RANKING order="8" place="8" resultid="3232" />
                    <RANKING order="9" place="-1" resultid="3894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1473" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6551" />
                    <RANKING order="2" place="2" resultid="4334" />
                    <RANKING order="3" place="3" resultid="1939" />
                    <RANKING order="4" place="4" resultid="3541" />
                    <RANKING order="5" place="5" resultid="2171" />
                    <RANKING order="6" place="6" resultid="3254" />
                    <RANKING order="7" place="7" resultid="2286" />
                    <RANKING order="8" place="-1" resultid="1871" />
                    <RANKING order="9" place="-1" resultid="2684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1474" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4804" />
                    <RANKING order="2" place="2" resultid="2532" />
                    <RANKING order="3" place="-1" resultid="3323" />
                    <RANKING order="4" place="-1" resultid="4034" />
                    <RANKING order="5" place="-1" resultid="4628" />
                    <RANKING order="6" place="-1" resultid="6035" />
                    <RANKING order="7" place="-1" resultid="1804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1475" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4363" />
                    <RANKING order="2" place="2" resultid="2716" />
                    <RANKING order="3" place="3" resultid="3771" />
                    <RANKING order="4" place="4" resultid="3965" />
                    <RANKING order="5" place="5" resultid="2108" />
                    <RANKING order="6" place="6" resultid="2920" />
                    <RANKING order="7" place="-1" resultid="1860" />
                    <RANKING order="8" place="-1" resultid="1834" />
                    <RANKING order="9" place="-1" resultid="3153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1476" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4590" />
                    <RANKING order="2" place="2" resultid="6023" />
                    <RANKING order="3" place="3" resultid="2516" />
                    <RANKING order="4" place="4" resultid="1954" />
                    <RANKING order="5" place="5" resultid="3816" />
                    <RANKING order="6" place="6" resultid="3216" />
                    <RANKING order="7" place="7" resultid="3913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1477" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2638" />
                    <RANKING order="2" place="2" resultid="2234" />
                    <RANKING order="3" place="-1" resultid="3944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1478" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1984" />
                    <RANKING order="2" place="2" resultid="3208" />
                    <RANKING order="3" place="3" resultid="3856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1479" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1480" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1481" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6299" daytime="20:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6300" daytime="20:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6301" daytime="20:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6302" daytime="20:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6303" daytime="20:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6304" daytime="20:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6305" daytime="20:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6306" daytime="20:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6307" daytime="20:40" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6308" daytime="20:45" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6309" daytime="20:45" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6310" daytime="20:50" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6311" daytime="20:50" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2012-11-25" daytime="09:00" name="Blok IV" number="4" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1483" daytime="09:00" gender="F" number="30" order="36" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1484" agemax="24" agemin="20" name="0: 20 - 24 lat" />
                <AGEGROUP agegroupid="1485" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3656" />
                    <RANKING order="2" place="2" resultid="4043" />
                    <RANKING order="3" place="3" resultid="4089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1486" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2859" />
                    <RANKING order="2" place="2" resultid="2392" />
                    <RANKING order="3" place="3" resultid="3481" />
                    <RANKING order="4" place="4" resultid="4059" />
                    <RANKING order="5" place="-1" resultid="4687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1487" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1488" agemax="44" agemin="40" name="D: 40 - 44 lat" />
                <AGEGROUP agegroupid="1489" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2140" />
                    <RANKING order="2" place="2" resultid="2563" />
                    <RANKING order="3" place="-1" resultid="3804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1490" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3781" />
                    <RANKING order="2" place="2" resultid="3621" />
                    <RANKING order="3" place="3" resultid="2003" />
                    <RANKING order="4" place="4" resultid="1961" />
                    <RANKING order="5" place="5" resultid="3468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1491" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2223" />
                    <RANKING order="2" place="2" resultid="1976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1492" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1878" />
                    <RANKING order="2" place="2" resultid="1969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1493" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1494" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1495" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1496" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1497" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6312" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6313" daytime="09:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6314" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6315" daytime="09:05" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1498" daytime="09:10" gender="M" number="31" order="37" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1499" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2755" />
                    <RANKING order="2" place="2" resultid="2021" />
                    <RANKING order="3" place="3" resultid="2078" />
                    <RANKING order="4" place="4" resultid="2803" />
                    <RANKING order="5" place="5" resultid="4616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1500" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3102" />
                    <RANKING order="2" place="2" resultid="3112" />
                    <RANKING order="3" place="3" resultid="4637" />
                    <RANKING order="4" place="4" resultid="2456" />
                    <RANKING order="5" place="5" resultid="2086" />
                    <RANKING order="6" place="6" resultid="2664" />
                    <RANKING order="7" place="7" resultid="4097" />
                    <RANKING order="8" place="-1" resultid="2668" />
                    <RANKING order="9" place="-1" resultid="3789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1501" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3486" />
                    <RANKING order="2" place="2" resultid="1787" />
                    <RANKING order="3" place="3" resultid="3643" />
                    <RANKING order="4" place="4" resultid="4715" />
                    <RANKING order="5" place="5" resultid="3369" />
                    <RANKING order="6" place="6" resultid="3649" />
                    <RANKING order="7" place="7" resultid="4077" />
                    <RANKING order="8" place="8" resultid="2509" />
                    <RANKING order="9" place="9" resultid="3238" />
                    <RANKING order="10" place="-1" resultid="3407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1502" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2494" />
                    <RANKING order="2" place="2" resultid="4027" />
                    <RANKING order="3" place="3" resultid="3562" />
                    <RANKING order="4" place="4" resultid="3182" />
                    <RANKING order="5" place="-1" resultid="2579" />
                    <RANKING order="6" place="-1" resultid="2852" />
                    <RANKING order="7" place="-1" resultid="4320" />
                    <RANKING order="8" place="-1" resultid="4608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1503" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2184" />
                    <RANKING order="2" place="2" resultid="3130" />
                    <RANKING order="3" place="3" resultid="4234" />
                    <RANKING order="4" place="4" resultid="3124" />
                    <RANKING order="5" place="-1" resultid="3895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1504" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1940" />
                    <RANKING order="2" place="2" resultid="4377" />
                    <RANKING order="3" place="3" resultid="2571" />
                    <RANKING order="4" place="4" resultid="3542" />
                    <RANKING order="5" place="5" resultid="2406" />
                    <RANKING order="6" place="6" resultid="1872" />
                    <RANKING order="7" place="-1" resultid="2677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1505" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4805" />
                    <RANKING order="2" place="2" resultid="3497" />
                    <RANKING order="3" place="3" resultid="2249" />
                    <RANKING order="4" place="4" resultid="2533" />
                    <RANKING order="5" place="5" resultid="1805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1506" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1861" />
                    <RANKING order="2" place="2" resultid="3225" />
                    <RANKING order="3" place="3" resultid="3849" />
                    <RANKING order="4" place="4" resultid="3738" />
                    <RANKING order="5" place="5" resultid="2921" />
                    <RANKING order="6" place="6" resultid="2910" />
                    <RANKING order="7" place="-1" resultid="1835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1507" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4675" />
                    <RANKING order="2" place="2" resultid="3586" />
                    <RANKING order="3" place="3" resultid="3914" />
                    <RANKING order="4" place="4" resultid="3217" />
                    <RANKING order="5" place="-1" resultid="3573" />
                    <RANKING order="6" place="-1" resultid="4591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1508" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2639" />
                    <RANKING order="2" place="2" resultid="1853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1509" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3161" />
                    <RANKING order="2" place="2" resultid="3209" />
                    <RANKING order="3" place="3" resultid="3857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1510" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1932" />
                    <RANKING order="2" place="2" resultid="4295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1511" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1512" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6316" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6317" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6318" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6319" daytime="09:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6320" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6321" daytime="09:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6322" daytime="09:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6323" daytime="09:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6324" daytime="09:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6325" daytime="09:30" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6326" daytime="09:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6327" daytime="09:30" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1513" daytime="09:35" gender="F" number="32" order="38" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1514" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2102" />
                    <RANKING order="2" place="2" resultid="2649" />
                    <RANKING order="3" place="3" resultid="3926" />
                    <RANKING order="4" place="4" resultid="2451" />
                    <RANKING order="5" place="5" resultid="2030" />
                    <RANKING order="6" place="6" resultid="2306" />
                    <RANKING order="7" place="7" resultid="3289" />
                    <RANKING order="8" place="8" resultid="2708" />
                    <RANKING order="9" place="-1" resultid="4738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1515" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3315" />
                    <RANKING order="2" place="2" resultid="3519" />
                    <RANKING order="3" place="3" resultid="1925" />
                    <RANKING order="4" place="4" resultid="4090" />
                    <RANKING order="5" place="5" resultid="4020" />
                    <RANKING order="6" place="6" resultid="4694" />
                    <RANKING order="7" place="7" resultid="2701" />
                    <RANKING order="8" place="-1" resultid="2891" />
                    <RANKING order="9" place="-1" resultid="4429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1516" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2860" />
                    <RANKING order="2" place="2" resultid="2828" />
                    <RANKING order="3" place="-1" resultid="4601" />
                    <RANKING order="4" place="-1" resultid="4688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4239" />
                    <RANKING order="2" place="2" resultid="3528" />
                    <RANKING order="3" place="3" resultid="3614" />
                    <RANKING order="4" place="4" resultid="4051" />
                    <RANKING order="5" place="5" resultid="3269" />
                    <RANKING order="6" place="6" resultid="2152" />
                    <RANKING order="7" place="7" resultid="3050" />
                    <RANKING order="8" place="-1" resultid="2841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1518" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4482" />
                    <RANKING order="2" place="2" resultid="4415" />
                    <RANKING order="3" place="3" resultid="4212" />
                    <RANKING order="4" place="4" resultid="4115" />
                    <RANKING order="5" place="5" resultid="3262" />
                    <RANKING order="6" place="6" resultid="2127" />
                    <RANKING order="7" place="7" resultid="2871" />
                    <RANKING order="8" place="-1" resultid="2884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1519" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2134" />
                    <RANKING order="2" place="2" resultid="4797" />
                    <RANKING order="3" place="3" resultid="2564" />
                    <RANKING order="4" place="4" resultid="4384" />
                    <RANKING order="5" place="5" resultid="2312" />
                    <RANKING order="6" place="6" resultid="4583" />
                    <RANKING order="7" place="7" resultid="4668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1520" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1847" />
                    <RANKING order="2" place="2" resultid="1841" />
                    <RANKING order="3" place="3" resultid="2004" />
                    <RANKING order="4" place="4" resultid="1772" />
                    <RANKING order="5" place="5" resultid="3475" />
                    <RANKING order="6" place="6" resultid="2819" />
                    <RANKING order="7" place="7" resultid="2998" />
                    <RANKING order="8" place="-1" resultid="3782" />
                    <RANKING order="9" place="-1" resultid="2740" />
                    <RANKING order="10" place="-1" resultid="1948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1521" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1825" />
                    <RANKING order="2" place="2" resultid="4149" />
                    <RANKING order="3" place="3" resultid="3138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1522" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4169" />
                    <RANKING order="2" place="2" resultid="2773" />
                    <RANKING order="3" place="3" resultid="3933" />
                    <RANKING order="4" place="4" resultid="4192" />
                    <RANKING order="5" place="5" resultid="2957" />
                    <RANKING order="6" place="6" resultid="1879" />
                    <RANKING order="7" place="7" resultid="4440" />
                    <RANKING order="8" place="8" resultid="2942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1523" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4174" />
                    <RANKING order="2" place="2" resultid="2164" />
                    <RANKING order="3" place="3" resultid="2949" />
                    <RANKING order="4" place="4" resultid="2935" />
                    <RANKING order="5" place="5" resultid="2964" />
                    <RANKING order="6" place="-1" resultid="4460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1524" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1525" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1526" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1527" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6328" daytime="09:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6329" daytime="09:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6330" daytime="09:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6331" daytime="09:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6332" daytime="09:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6333" daytime="09:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6334" daytime="09:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6335" daytime="09:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6336" daytime="09:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6337" daytime="09:45" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6338" daytime="09:45" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6339" daytime="09:45" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6340" daytime="09:50" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1528" daytime="09:50" gender="M" number="33" order="39" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1529" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3877" />
                    <RANKING order="2" place="2" resultid="2022" />
                    <RANKING order="3" place="3" resultid="3066" />
                    <RANKING order="4" place="4" resultid="2804" />
                    <RANKING order="5" place="5" resultid="2419" />
                    <RANKING order="6" place="6" resultid="2215" />
                    <RANKING order="7" place="7" resultid="4622" />
                    <RANKING order="8" place="8" resultid="2657" />
                    <RANKING order="9" place="-1" resultid="4532" />
                    <RANKING order="10" place="-1" resultid="4547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1530" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2727" />
                    <RANKING order="2" place="2" resultid="3880" />
                    <RANKING order="3" place="3" resultid="4315" />
                    <RANKING order="4" place="4" resultid="4701" />
                    <RANKING order="5" place="5" resultid="3862" />
                    <RANKING order="6" place="6" resultid="3400" />
                    <RANKING order="7" place="7" resultid="3415" />
                    <RANKING order="8" place="8" resultid="2117" />
                    <RANKING order="9" place="9" resultid="4108" />
                    <RANKING order="10" place="10" resultid="2586" />
                    <RANKING order="11" place="11" resultid="4098" />
                    <RANKING order="12" place="-1" resultid="3072" />
                    <RANKING order="13" place="-1" resultid="3104" />
                    <RANKING order="14" place="-1" resultid="3462" />
                    <RANKING order="15" place="-1" resultid="3790" />
                    <RANKING order="16" place="-1" resultid="4435" />
                    <RANKING order="17" place="-1" resultid="4541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1531" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4445" />
                    <RANKING order="2" place="2" resultid="4711" />
                    <RANKING order="3" place="3" resultid="4102" />
                    <RANKING order="4" place="4" resultid="4345" />
                    <RANKING order="5" place="5" resultid="3487" />
                    <RANKING order="6" place="6" resultid="3095" />
                    <RANKING order="7" place="7" resultid="3370" />
                    <RANKING order="8" place="8" resultid="4767" />
                    <RANKING order="9" place="9" resultid="2308" />
                    <RANKING order="10" place="10" resultid="3350" />
                    <RANKING order="11" place="11" resultid="3106" />
                    <RANKING order="12" place="12" resultid="4469" />
                    <RANKING order="13" place="13" resultid="3580" />
                    <RANKING order="14" place="14" resultid="3823" />
                    <RANKING order="15" place="15" resultid="3380" />
                    <RANKING order="16" place="16" resultid="3567" />
                    <RANKING order="17" place="17" resultid="4357" />
                    <RANKING order="18" place="18" resultid="3375" />
                    <RANKING order="19" place="19" resultid="3239" />
                    <RANKING order="20" place="20" resultid="2254" />
                    <RANKING order="21" place="21" resultid="3921" />
                    <RANKING order="22" place="-1" resultid="4810" />
                    <RANKING order="23" place="-1" resultid="3359" />
                    <RANKING order="24" place="-1" resultid="3098" />
                    <RANKING order="25" place="-1" resultid="3292" />
                    <RANKING order="26" place="-1" resultid="3354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1532" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3490" />
                    <RANKING order="2" place="2" resultid="4817" />
                    <RANKING order="3" place="3" resultid="2486" />
                    <RANKING order="4" place="4" resultid="4028" />
                    <RANKING order="5" place="5" resultid="3306" />
                    <RANKING order="6" place="6" resultid="3387" />
                    <RANKING order="7" place="7" resultid="4397" />
                    <RANKING order="8" place="8" resultid="3563" />
                    <RANKING order="9" place="9" resultid="3116" />
                    <RANKING order="10" place="10" resultid="2398" />
                    <RANKING order="11" place="11" resultid="2439" />
                    <RANKING order="12" place="12" resultid="2914" />
                    <RANKING order="13" place="13" resultid="2837" />
                    <RANKING order="14" place="14" resultid="4609" />
                    <RANKING order="15" place="15" resultid="3493" />
                    <RANKING order="16" place="16" resultid="1778" />
                    <RANKING order="17" place="-1" resultid="2299" />
                    <RANKING order="18" place="-1" resultid="2466" />
                    <RANKING order="19" place="-1" resultid="3983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1533" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2825" />
                    <RANKING order="2" place="2" resultid="2780" />
                    <RANKING order="3" place="3" resultid="1754" />
                    <RANKING order="4" place="4" resultid="2192" />
                    <RANKING order="5" place="5" resultid="3131" />
                    <RANKING order="6" place="6" resultid="3170" />
                    <RANKING order="7" place="7" resultid="2479" />
                    <RANKING order="8" place="8" resultid="2525" />
                    <RANKING order="9" place="9" resultid="2730" />
                    <RANKING order="10" place="10" resultid="3896" />
                    <RANKING order="11" place="11" resultid="3233" />
                    <RANKING order="12" place="12" resultid="2045" />
                    <RANKING order="13" place="13" resultid="3977" />
                    <RANKING order="14" place="14" resultid="3247" />
                    <RANKING order="15" place="-1" resultid="4328" />
                    <RANKING order="16" place="-1" resultid="1746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1534" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3509" />
                    <RANKING order="2" place="2" resultid="3549" />
                    <RANKING order="3" place="3" resultid="2685" />
                    <RANKING order="4" place="4" resultid="2785" />
                    <RANKING order="5" place="5" resultid="1941" />
                    <RANKING order="6" place="6" resultid="4335" />
                    <RANKING order="7" place="7" resultid="4661" />
                    <RANKING order="8" place="8" resultid="2430" />
                    <RANKING order="9" place="9" resultid="3255" />
                    <RANKING order="10" place="10" resultid="2172" />
                    <RANKING order="11" place="11" resultid="2267" />
                    <RANKING order="12" place="12" resultid="2274" />
                    <RANKING order="13" place="13" resultid="3716" />
                    <RANKING order="14" place="14" resultid="4342" />
                    <RANKING order="15" place="-1" resultid="4083" />
                    <RANKING order="16" place="-1" resultid="2384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1535" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4309" />
                    <RANKING order="2" place="2" resultid="2435" />
                    <RANKING order="3" place="3" resultid="3810" />
                    <RANKING order="4" place="4" resultid="4719" />
                    <RANKING order="5" place="5" resultid="2903" />
                    <RANKING order="6" place="6" resultid="1884" />
                    <RANKING order="7" place="7" resultid="4629" />
                    <RANKING order="8" place="8" resultid="2539" />
                    <RANKING order="9" place="9" resultid="6036" />
                    <RANKING order="10" place="-1" resultid="2835" />
                    <RANKING order="11" place="-1" resultid="3324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1536" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1797" />
                    <RANKING order="2" place="2" resultid="2767" />
                    <RANKING order="3" place="3" resultid="2061" />
                    <RANKING order="4" place="4" resultid="4144" />
                    <RANKING order="5" place="5" resultid="2109" />
                    <RANKING order="6" place="6" resultid="3005" />
                    <RANKING order="7" place="-1" resultid="4070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1537" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3722" />
                    <RANKING order="2" place="2" resultid="3587" />
                    <RANKING order="3" place="3" resultid="4676" />
                    <RANKING order="4" place="4" resultid="4163" />
                    <RANKING order="5" place="5" resultid="2124" />
                    <RANKING order="6" place="6" resultid="4351" />
                    <RANKING order="7" place="7" resultid="4218" />
                    <RANKING order="8" place="8" resultid="2621" />
                    <RANKING order="9" place="-1" resultid="4224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1538" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2640" />
                    <RANKING order="2" place="2" resultid="2235" />
                    <RANKING order="3" place="3" resultid="1854" />
                    <RANKING order="4" place="4" resultid="2202" />
                    <RANKING order="5" place="5" resultid="2206" />
                    <RANKING order="6" place="6" resultid="2816" />
                    <RANKING order="7" place="-1" resultid="2977" />
                    <RANKING order="8" place="-1" resultid="4371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1539" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4160" />
                    <RANKING order="2" place="2" resultid="1985" />
                    <RANKING order="3" place="3" resultid="3601" />
                    <RANKING order="4" place="4" resultid="3201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1540" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3701" />
                    <RANKING order="2" place="2" resultid="4724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1541" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3766" />
                    <RANKING order="2" place="2" resultid="1667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1542" agemax="-1" agemin="85" name="M: 85 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1866" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6341" daytime="09:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6342" daytime="09:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6343" daytime="09:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6344" daytime="09:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6345" daytime="09:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6346" daytime="09:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6347" daytime="10:00" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6348" daytime="10:00" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6349" daytime="10:00" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6350" daytime="10:00" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6351" daytime="10:00" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6352" daytime="10:05" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6353" daytime="10:05" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6354" daytime="10:05" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="6355" daytime="10:05" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="6356" daytime="10:05" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="6357" daytime="10:10" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="6358" daytime="10:10" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="6359" daytime="10:10" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="6360" daytime="10:10" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="6361" daytime="10:10" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="6362" daytime="10:10" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="6363" daytime="10:15" number="23" order="23" status="OFFICIAL" />
                <HEAT heatid="6364" daytime="10:15" number="24" order="24" status="OFFICIAL" />
                <HEAT heatid="6365" daytime="10:15" number="25" order="25" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1543" daytime="10:15" gender="F" number="34" order="40" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1544" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2452" />
                    <RANKING order="2" place="2" resultid="2709" />
                    <RANKING order="3" place="3" resultid="3629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1545" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2242" />
                    <RANKING order="2" place="2" resultid="4044" />
                    <RANKING order="3" place="3" resultid="4695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1546" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3636" />
                    <RANKING order="2" place="2" resultid="2393" />
                    <RANKING order="3" place="3" resultid="4602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1547" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3999" />
                    <RANKING order="2" place="2" resultid="2794" />
                    <RANKING order="3" place="3" resultid="4052" />
                    <RANKING order="4" place="-1" resultid="4303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1548" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4213" />
                    <RANKING order="2" place="2" resultid="2296" />
                    <RANKING order="3" place="3" resultid="4116" />
                    <RANKING order="4" place="4" resultid="3299" />
                    <RANKING order="5" place="-1" resultid="2264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1549" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2135" />
                    <RANKING order="2" place="2" resultid="2414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1550" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3840" />
                    <RANKING order="2" place="2" resultid="1842" />
                    <RANKING order="3" place="3" resultid="1993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1551" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4150" />
                    <RANKING order="2" place="2" resultid="2927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1552" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4170" />
                    <RANKING order="2" place="2" resultid="2943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1553" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1554" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4643" />
                    <RANKING order="2" place="2" resultid="1817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1555" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1556" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1557" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6366" daytime="10:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6367" daytime="10:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6368" daytime="10:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6369" daytime="10:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6370" daytime="10:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6371" daytime="10:40" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1558" daytime="10:45" gender="M" number="35" order="41" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1559" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2756" />
                    <RANKING order="2" place="2" resultid="4617" />
                    <RANKING order="3" place="3" resultid="4548" />
                    <RANKING order="4" place="-1" resultid="1737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1560" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3113" />
                    <RANKING order="2" place="2" resultid="2631" />
                    <RANKING order="3" place="3" resultid="3278" />
                    <RANKING order="4" place="-1" resultid="2736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1561" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3287" />
                    <RANKING order="2" place="2" resultid="3644" />
                    <RANKING order="3" place="3" resultid="3608" />
                    <RANKING order="4" place="4" resultid="3408" />
                    <RANKING order="5" place="5" resultid="3341" />
                    <RANKING order="6" place="-1" resultid="3333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1562" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2487" />
                    <RANKING order="2" place="2" resultid="4398" />
                    <RANKING order="3" place="3" resultid="2555" />
                    <RANKING order="4" place="-1" resultid="4321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1563" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4206" />
                    <RANKING order="2" place="2" resultid="2053" />
                    <RANKING order="3" place="3" resultid="3016" />
                    <RANKING order="4" place="4" resultid="2526" />
                    <RANKING order="5" place="5" resultid="3831" />
                    <RANKING order="6" place="6" resultid="1765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1564" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4336" />
                    <RANKING order="2" place="2" resultid="4662" />
                    <RANKING order="3" place="3" resultid="2686" />
                    <RANKING order="4" place="4" resultid="2431" />
                    <RANKING order="5" place="5" resultid="2572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1565" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4035" />
                    <RANKING order="2" place="2" resultid="3729" />
                    <RANKING order="3" place="3" resultid="2095" />
                    <RANKING order="4" place="4" resultid="2534" />
                    <RANKING order="5" place="5" resultid="3043" />
                    <RANKING order="6" place="6" resultid="6037" />
                    <RANKING order="7" place="7" resultid="4408" />
                    <RANKING order="8" place="-1" resultid="4008" />
                    <RANKING order="9" place="-1" resultid="2250" />
                    <RANKING order="10" place="-1" resultid="2069" />
                    <RANKING order="11" place="-1" resultid="2904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1566" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4364" />
                    <RANKING order="2" place="2" resultid="3772" />
                    <RANKING order="3" place="3" resultid="3966" />
                    <RANKING order="4" place="4" resultid="3535" />
                    <RANKING order="5" place="5" resultid="3739" />
                    <RANKING order="6" place="6" resultid="3226" />
                    <RANKING order="7" place="7" resultid="2110" />
                    <RANKING order="8" place="-1" resultid="3154" />
                    <RANKING order="9" place="-1" resultid="2717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1567" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4476" />
                    <RANKING order="2" place="2" resultid="3723" />
                    <RANKING order="3" place="3" resultid="2517" />
                    <RANKING order="4" place="4" resultid="3915" />
                    <RANKING order="5" place="5" resultid="3817" />
                    <RANKING order="6" place="6" resultid="3012" />
                    <RANKING order="7" place="7" resultid="6544" />
                    <RANKING order="8" place="-1" resultid="3958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1568" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3952" />
                    <RANKING order="2" place="2" resultid="4187" />
                    <RANKING order="3" place="3" resultid="3945" />
                    <RANKING order="4" place="4" resultid="2991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1569" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3210" />
                    <RANKING order="2" place="2" resultid="3602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1570" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1571" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1572" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6372" daytime="10:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6373" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6374" daytime="10:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6375" daytime="11:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6376" daytime="11:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6377" daytime="11:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6378" daytime="11:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6379" daytime="11:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6380" daytime="11:20" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6381" daytime="11:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6382" daytime="11:25" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1588" daytime="11:30" gender="X" number="36" order="42" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1589" agemax="119" agemin="100" name="A: 100 - 119 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="1590" agemax="159" agemin="120" name="B: 120 - 159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3668" />
                    <RANKING order="2" place="2" resultid="2323" />
                    <RANKING order="3" place="3" resultid="4494" />
                    <RANKING order="4" place="4" resultid="4122" />
                    <RANKING order="5" place="5" resultid="3501" />
                    <RANKING order="6" place="6" resultid="4124" />
                    <RANKING order="7" place="7" resultid="4733" />
                    <RANKING order="8" place="8" resultid="4495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1591" agemax="199" agemin="160" name="C: 160 - 199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2324" />
                    <RANKING order="2" place="2" resultid="4261" />
                    <RANKING order="3" place="3" resultid="4493" />
                    <RANKING order="4" place="4" resultid="3272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1592" agemax="239" agemin="200" name="D: 200 - 239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2325" />
                    <RANKING order="2" place="2" resultid="1895" />
                    <RANKING order="3" place="3" resultid="3022" />
                    <RANKING order="4" place="4" resultid="3164" />
                    <RANKING order="5" place="-1" resultid="2326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1593" agemax="279" agemin="240" name="E: 240 - 279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="4734" />
                    <RANKING order="3" place="3" resultid="1890" />
                    <RANKING order="4" place="4" resultid="1722" />
                    <RANKING order="5" place="5" resultid="2327" />
                    <RANKING order="6" place="6" resultid="3023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1594" agemax="-1" agemin="280" name="F: 280 lat i starsi" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4259" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6535" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6536" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6537" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6538" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1595" daytime="11:40" gender="F" number="37" order="43" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1596" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2103" />
                    <RANKING order="2" place="2" resultid="2723" />
                    <RANKING order="3" place="3" resultid="6501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1597" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3316" />
                    <RANKING order="2" place="2" resultid="3657" />
                    <RANKING order="3" place="3" resultid="2280" />
                    <RANKING order="4" place="4" resultid="4430" />
                    <RANKING order="5" place="5" resultid="2210" />
                    <RANKING order="6" place="6" resultid="4575" />
                    <RANKING order="7" place="-1" resultid="2892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1598" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4064" />
                    <RANKING order="2" place="2" resultid="2039" />
                    <RANKING order="3" place="3" resultid="3515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3615" />
                    <RANKING order="2" place="2" resultid="3529" />
                    <RANKING order="3" place="3" resultid="3270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4199" />
                    <RANKING order="2" place="2" resultid="3263" />
                    <RANKING order="3" place="3" resultid="2265" />
                    <RANKING order="4" place="-1" resultid="2885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4385" />
                    <RANKING order="2" place="2" resultid="4584" />
                    <RANKING order="3" place="3" resultid="4455" />
                    <RANKING order="4" place="4" resultid="4669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2144" />
                    <RANKING order="2" place="2" resultid="1848" />
                    <RANKING order="3" place="3" resultid="4681" />
                    <RANKING order="4" place="4" resultid="1773" />
                    <RANKING order="5" place="5" resultid="3469" />
                    <RANKING order="6" place="6" resultid="2999" />
                    <RANKING order="7" place="7" resultid="3146" />
                    <RANKING order="8" place="-1" resultid="3622" />
                    <RANKING order="9" place="-1" resultid="4230" />
                    <RANKING order="10" place="-1" resultid="1962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3939" />
                    <RANKING order="2" place="2" resultid="1977" />
                    <RANKING order="3" place="3" resultid="3139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3934" />
                    <RANKING order="2" place="2" resultid="2158" />
                    <RANKING order="3" place="3" resultid="1970" />
                    <RANKING order="4" place="4" resultid="2810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4154" />
                    <RANKING order="2" place="2" resultid="4179" />
                    <RANKING order="3" place="3" resultid="2165" />
                    <RANKING order="4" place="4" resultid="2936" />
                    <RANKING order="5" place="5" resultid="2965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1606" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1818" />
                    <RANKING order="2" place="2" resultid="2971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1607" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1608" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1609" agemax="-1" agemin="85" name="M: 85 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1980" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6502" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6503" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6504" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6505" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6506" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6507" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6508" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6509" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6510" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1610" daytime="12:00" gender="M" number="38" order="44" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1611" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4566" />
                    <RANKING order="2" place="2" resultid="4536" />
                    <RANKING order="3" place="3" resultid="3067" />
                    <RANKING order="4" place="-1" resultid="1738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1612" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4558" />
                    <RANKING order="2" place="2" resultid="4466" />
                    <RANKING order="3" place="3" resultid="2653" />
                    <RANKING order="4" place="4" resultid="2118" />
                    <RANKING order="5" place="5" resultid="3279" />
                    <RANKING order="6" place="6" resultid="3416" />
                    <RANKING order="7" place="7" resultid="3394" />
                    <RANKING order="8" place="8" resultid="3401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1613" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6571" />
                    <RANKING order="2" place="2" resultid="3364" />
                    <RANKING order="3" place="3" resultid="1791" />
                    <RANKING order="4" place="4" resultid="2510" />
                    <RANKING order="5" place="5" resultid="3581" />
                    <RANKING order="6" place="6" resultid="3342" />
                    <RANKING order="7" place="7" resultid="3346" />
                    <RANKING order="8" place="-1" resultid="4078" />
                    <RANKING order="9" place="-1" resultid="3240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1614" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2580" />
                    <RANKING order="2" place="2" resultid="2547" />
                    <RANKING order="3" place="3" resultid="4818" />
                    <RANKING order="4" place="4" resultid="2317" />
                    <RANKING order="5" place="5" resultid="2502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1615" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3452" />
                    <RANKING order="2" place="2" resultid="4013" />
                    <RANKING order="3" place="3" resultid="2228" />
                    <RANKING order="4" place="4" resultid="3017" />
                    <RANKING order="5" place="5" resultid="3125" />
                    <RANKING order="6" place="6" resultid="3832" />
                    <RANKING order="7" place="7" resultid="3248" />
                    <RANKING order="8" place="8" resultid="2444" />
                    <RANKING order="9" place="9" resultid="3978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1616" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3510" />
                    <RANKING order="2" place="2" resultid="3972" />
                    <RANKING order="3" place="3" resultid="3543" />
                    <RANKING order="4" place="4" resultid="2268" />
                    <RANKING order="5" place="5" resultid="2173" />
                    <RANKING order="6" place="6" resultid="4343" />
                    <RANKING order="7" place="7" resultid="3256" />
                    <RANKING order="8" place="8" resultid="1873" />
                    <RANKING order="9" place="-1" resultid="2385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1617" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4036" />
                    <RANKING order="2" place="2" resultid="3554" />
                    <RANKING order="3" place="3" resultid="2540" />
                    <RANKING order="4" place="4" resultid="1885" />
                    <RANKING order="5" place="5" resultid="2180" />
                    <RANKING order="6" place="-1" resultid="4630" />
                    <RANKING order="7" place="-1" resultid="4310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1618" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2747" />
                    <RANKING order="2" place="2" resultid="2832" />
                    <RANKING order="3" place="3" resultid="2768" />
                    <RANKING order="4" place="4" resultid="1836" />
                    <RANKING order="5" place="5" resultid="3661" />
                    <RANKING order="6" place="6" resultid="3732" />
                    <RANKING order="7" place="7" resultid="3006" />
                    <RANKING order="8" place="8" resultid="2922" />
                    <RANKING order="9" place="9" resultid="3058" />
                    <RANKING order="10" place="10" resultid="3155" />
                    <RANKING order="11" place="-1" resultid="1798" />
                    <RANKING order="12" place="-1" resultid="4071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1619" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4592" />
                    <RANKING order="2" place="2" resultid="1829" />
                    <RANKING order="3" place="3" resultid="1955" />
                    <RANKING order="4" place="4" resultid="3818" />
                    <RANKING order="5" place="5" resultid="2303" />
                    <RANKING order="6" place="-1" resultid="3574" />
                    <RANKING order="7" place="-1" resultid="4242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1620" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3953" />
                    <RANKING order="2" place="2" resultid="2690" />
                    <RANKING order="3" place="3" resultid="2992" />
                    <RANKING order="4" place="4" resultid="2817" />
                    <RANKING order="5" place="-1" resultid="2978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1621" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4161" />
                    <RANKING order="2" place="2" resultid="4183" />
                    <RANKING order="3" place="3" resultid="1986" />
                    <RANKING order="4" place="4" resultid="3162" />
                    <RANKING order="5" place="5" resultid="3202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1622" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4296" />
                    <RANKING order="2" place="2" resultid="4725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1623" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1624" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6395" daytime="12:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6396" daytime="12:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6397" daytime="12:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6398" daytime="12:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6399" daytime="12:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6400" daytime="12:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6401" daytime="12:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6402" daytime="12:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6403" daytime="12:20" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6404" daytime="12:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6405" daytime="12:25" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6406" daytime="12:25" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6407" daytime="12:30" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6408" daytime="12:30" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1625" daytime="12:30" gender="F" number="39" order="45" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1626" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2031" />
                    <RANKING order="2" place="2" resultid="3927" />
                    <RANKING order="3" place="3" resultid="3630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1627" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2243" />
                    <RANKING order="2" place="2" resultid="4576" />
                    <RANKING order="3" place="3" resultid="4423" />
                    <RANKING order="4" place="4" resultid="2702" />
                    <RANKING order="5" place="-1" resultid="4021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1628" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2040" />
                    <RANKING order="2" place="2" resultid="4060" />
                    <RANKING order="3" place="3" resultid="3482" />
                    <RANKING order="4" place="4" resultid="4450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1629" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1659" />
                    <RANKING order="2" place="2" resultid="3051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1630" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4200" />
                    <RANKING order="2" place="2" resultid="4416" />
                    <RANKING order="3" place="3" resultid="2297" />
                    <RANKING order="4" place="4" resultid="3300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1631" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2471" />
                    <RANKING order="2" place="2" resultid="4798" />
                    <RANKING order="3" place="3" resultid="2415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1632" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3841" />
                    <RANKING order="2" place="2" resultid="1949" />
                    <RANKING order="3" place="3" resultid="1994" />
                    <RANKING order="4" place="4" resultid="2820" />
                    <RANKING order="5" place="5" resultid="3147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2224" />
                    <RANKING order="2" place="2" resultid="2928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2958" />
                    <RANKING order="2" place="2" resultid="4441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="69" agemin="65" name="I: 65 - 69 lat" />
                <AGEGROUP agegroupid="1636" agemax="74" agemin="70" name="J: 70 - 74 lat" />
                <AGEGROUP agegroupid="1637" agemax="79" agemin="75" name="K: 75 - 79 lat" />
                <AGEGROUP agegroupid="1638" agemax="84" agemin="80" name="L: 80 - 84 lat" />
                <AGEGROUP agegroupid="1639" agemax="-1" agemin="85" name="M: 85 lat i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6554" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6555" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6556" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6557" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6558" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1640" daytime="13:15" gender="M" number="40" order="46" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1641" agemax="24" agemin="20" name="0: 20 - 24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3878" />
                    <RANKING order="2" place="2" resultid="4567" />
                    <RANKING order="3" place="3" resultid="2079" />
                    <RANKING order="4" place="4" resultid="2420" />
                    <RANKING order="5" place="5" resultid="2216" />
                    <RANKING order="6" place="-1" resultid="4552" />
                    <RANKING order="7" place="-1" resultid="4704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1642" agemax="29" agemin="25" name="A: 25 - 25 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4638" />
                    <RANKING order="2" place="2" resultid="2087" />
                    <RANKING order="3" place="3" resultid="3906" />
                    <RANKING order="4" place="4" resultid="3863" />
                    <RANKING order="5" place="-1" resultid="2425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1643" agemax="34" agemin="30" name="B: 30 - 34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3334" />
                    <RANKING order="2" place="2" resultid="3824" />
                    <RANKING order="3" place="3" resultid="1783" />
                    <RANKING order="4" place="4" resultid="4358" />
                    <RANKING order="5" place="5" resultid="3650" />
                    <RANKING order="6" place="6" resultid="2188" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1644" agemax="39" agemin="35" name="C: 35 - 39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2495" />
                    <RANKING order="2" place="2" resultid="2467" />
                    <RANKING order="3" place="3" resultid="3307" />
                    <RANKING order="4" place="4" resultid="3388" />
                    <RANKING order="5" place="5" resultid="3117" />
                    <RANKING order="6" place="6" resultid="2556" />
                    <RANKING order="7" place="7" resultid="2399" />
                    <RANKING order="8" place="-1" resultid="2548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1645" agemax="44" agemin="40" name="D: 40 - 44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3453" />
                    <RANKING order="2" place="2" resultid="3171" />
                    <RANKING order="3" place="3" resultid="2480" />
                    <RANKING order="4" place="4" resultid="2054" />
                    <RANKING order="5" place="5" resultid="3866" />
                    <RANKING order="6" place="6" resultid="2046" />
                    <RANKING order="7" place="7" resultid="3234" />
                    <RANKING order="8" place="-1" resultid="1747" />
                    <RANKING order="9" place="-1" resultid="4329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1646" agemax="49" agemin="45" name="E: 45 - 49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4378" />
                    <RANKING order="2" place="2" resultid="3550" />
                    <RANKING order="3" place="3" resultid="2407" />
                    <RANKING order="4" place="4" resultid="2275" />
                    <RANKING order="5" place="5" resultid="2287" />
                    <RANKING order="6" place="-1" resultid="2696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1647" agemax="54" agemin="50" name="F: 50 - 54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2436" />
                    <RANKING order="2" place="2" resultid="6572" />
                    <RANKING order="3" place="3" resultid="1806" />
                    <RANKING order="4" place="4" resultid="2181" />
                    <RANKING order="5" place="5" resultid="4409" />
                    <RANKING order="6" place="-1" resultid="4806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1648" agemax="59" agemin="55" name="G: 55 - 59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2762" />
                    <RANKING order="2" place="2" resultid="3850" />
                    <RANKING order="3" place="3" resultid="2748" />
                    <RANKING order="4" place="4" resultid="4145" />
                    <RANKING order="5" place="5" resultid="2062" />
                    <RANKING order="6" place="6" resultid="3536" />
                    <RANKING order="7" place="7" resultid="3059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1649" agemax="64" agemin="60" name="H: 60 - 64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4477" />
                    <RANKING order="2" place="2" resultid="2518" />
                    <RANKING order="3" place="3" resultid="3959" />
                    <RANKING order="4" place="4" resultid="2125" />
                    <RANKING order="5" place="5" resultid="2984" />
                    <RANKING order="6" place="6" resultid="3218" />
                    <RANKING order="7" place="-1" resultid="6545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1650" agemax="69" agemin="65" name="I: 65 - 69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2236" />
                    <RANKING order="2" place="2" resultid="4372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1651" agemax="74" agemin="70" name="J: 70 - 74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1652" agemax="79" agemin="75" name="K: 75 - 79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1653" agemax="84" agemin="80" name="L: 80 - 84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2626" />
                    <RANKING order="2" place="2" resultid="1668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6517" agemax="89" agemin="85" name="M: 85 - 89 lat" />
                <AGEGROUP agegroupid="1654" agemax="-1" agemin="90" name="N: 90 lat i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1867" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6559" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6560" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6561" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6562" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6563" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6564" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6565" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6566" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6567" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6568" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6569" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6570" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" name="AZS Almamer" nation="POL">
          <CONTACT name="soltyk judyta" />
          <ATHLETES>
            <ATHLETE birthdate="1974-11-19" firstname="Judyta" gender="F" lastname="Sołtyk" nation="POL" athleteid="1656">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. C" eventid="1122" points="696" swimtime="00:10:32.00" resultid="1657" heatid="6445" lane="2" entrytime="00:10:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:13.80" />
                    <SPLIT distance="150" swimtime="00:01:52.56" />
                    <SPLIT distance="200" swimtime="00:02:32.10" />
                    <SPLIT distance="250" swimtime="00:03:11.99" />
                    <SPLIT distance="300" swimtime="00:03:51.98" />
                    <SPLIT distance="350" swimtime="00:04:32.06" />
                    <SPLIT distance="400" swimtime="00:05:12.72" />
                    <SPLIT distance="450" swimtime="00:05:53.12" />
                    <SPLIT distance="500" swimtime="00:06:33.59" />
                    <SPLIT distance="550" swimtime="00:07:13.94" />
                    <SPLIT distance="600" swimtime="00:07:54.12" />
                    <SPLIT distance="650" swimtime="00:08:34.44" />
                    <SPLIT distance="700" swimtime="00:09:14.58" />
                    <SPLIT distance="750" swimtime="00:09:54.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="617" reactiontime="+84" swimtime="00:02:27.78" resultid="1658" heatid="6277" lane="6" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:10.19" />
                    <SPLIT distance="150" swimtime="00:01:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="648" reactiontime="+84" swimtime="00:05:09.50" resultid="1659" heatid="6558" lane="5" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="150" swimtime="00:01:51.79" />
                    <SPLIT distance="200" swimtime="00:02:31.16" />
                    <SPLIT distance="250" swimtime="00:03:10.91" />
                    <SPLIT distance="300" swimtime="00:03:50.75" />
                    <SPLIT distance="350" swimtime="00:04:30.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="WOPR Kutno" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1932-01-01" firstname="Kazimierz" gender="M" lastname="From" nation="POL" athleteid="1661">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. L" eventid="1137" points="262" swimtime="00:22:38.64" resultid="1662" heatid="6447" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:32.60" />
                    <SPLIT distance="200" swimtime="00:05:25.09" />
                    <SPLIT distance="300" swimtime="00:08:22.82" />
                    <SPLIT distance="400" swimtime="00:11:15.22" />
                    <SPLIT distance="500" swimtime="00:16:06.89" />
                    <SPLIT distance="600" swimtime="00:17:00.62" />
                    <SPLIT distance="700" swimtime="00:19:53.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="162" reactiontime="+104" swimtime="00:01:15.14" resultid="1663" heatid="6126" lane="5" />
                <RESULT eventid="1272" points="206" reactiontime="+112" swimtime="00:02:10.99" resultid="1664" heatid="6159" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="167" reactiontime="+88" swimtime="00:02:48.68" resultid="1665" heatid="6249" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="262" reactiontime="+120" swimtime="00:05:00.84" resultid="1666" heatid="6278" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.47" />
                    <SPLIT distance="100" swimtime="00:02:25.69" />
                    <SPLIT distance="150" swimtime="00:03:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="201" reactiontime="+117" swimtime="00:00:56.54" resultid="1667" heatid="6341" lane="5" />
                <RESULT eventid="1640" points="248" reactiontime="+125" swimtime="00:10:55.37" resultid="1668" heatid="6559" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.79" />
                    <SPLIT distance="100" swimtime="00:02:17.57" />
                    <SPLIT distance="150" swimtime="00:03:37.82" />
                    <SPLIT distance="200" swimtime="00:05:02.82" />
                    <SPLIT distance="250" swimtime="00:06:31.85" />
                    <SPLIT distance="300" swimtime="00:08:01.58" />
                    <SPLIT distance="350" swimtime="00:09:32.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Gdynia Masters" nation="POL">
          <CONTACT email="misiek@am.gdynia.pl" name="Mysiak Katarzyna" />
          <ATHLETES>
            <ATHLETE birthdate="1961-01-01" firstname="Mysiak" gender="F" lastname="Katarzyna" nation="POL" athleteid="1943">
              <RESULTS>
                <RESULT eventid="1122" points="425" swimtime="00:13:57.84" resultid="1944" heatid="6443" lane="2" entrytime="00:14:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.22" />
                    <SPLIT distance="100" swimtime="00:01:36.60" />
                    <SPLIT distance="200" swimtime="00:03:22.50" />
                    <SPLIT distance="300" swimtime="00:05:09.61" />
                    <SPLIT distance="400" swimtime="00:06:56.66" />
                    <SPLIT distance="500" swimtime="00:08:43.65" />
                    <SPLIT distance="600" swimtime="00:10:30.55" />
                    <SPLIT distance="700" swimtime="00:12:16.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="469" reactiontime="+77" swimtime="00:00:44.51" resultid="1945" heatid="6122" lane="6" entrytime="00:00:44.00" />
                <RESULT eventid="1257" points="434" reactiontime="+98" swimtime="00:01:25.87" resultid="1946" heatid="6151" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="431" reactiontime="+114" swimtime="00:03:09.68" resultid="1947" heatid="6274" lane="4" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                    <SPLIT distance="100" swimtime="00:01:31.09" />
                    <SPLIT distance="150" swimtime="00:02:21.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="1948" heatid="6334" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1625" points="467" reactiontime="+105" swimtime="00:06:38.20" resultid="1949" heatid="6556" lane="6" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                    <SPLIT distance="100" swimtime="00:01:32.51" />
                    <SPLIT distance="150" swimtime="00:02:23.09" />
                    <SPLIT distance="200" swimtime="00:03:14.23" />
                    <SPLIT distance="250" swimtime="00:04:05.86" />
                    <SPLIT distance="300" swimtime="00:04:56.58" />
                    <SPLIT distance="350" swimtime="00:05:48.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Czeslaw" gender="M" lastname="Mikolajczyk" nation="POL" athleteid="1950">
              <RESULTS>
                <RESULT eventid="1092" points="471" reactiontime="+104" swimtime="00:07:27.43" resultid="1951" heatid="6487" lane="6" entrytime="00:07:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.97" />
                    <SPLIT distance="100" swimtime="00:01:48.21" />
                    <SPLIT distance="150" swimtime="00:02:47.61" />
                    <SPLIT distance="200" swimtime="00:03:45.79" />
                    <SPLIT distance="250" swimtime="00:05:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="532" reactiontime="+92" swimtime="00:03:37.76" resultid="1952" heatid="6110" lane="2" entrytime="00:03:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.51" />
                    <SPLIT distance="100" swimtime="00:01:43.68" />
                    <SPLIT distance="150" swimtime="00:02:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="439" reactiontime="+97" swimtime="00:00:45.07" resultid="1953" heatid="6207" lane="6" entrytime="00:00:44.00" />
                <RESULT eventid="1467" points="469" reactiontime="+94" swimtime="00:03:27.36" resultid="1954" heatid="6302" lane="6" entrytime="00:03:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                    <SPLIT distance="100" swimtime="00:01:45.04" />
                    <SPLIT distance="150" swimtime="00:02:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="485" reactiontime="+92" swimtime="00:01:40.49" resultid="1955" heatid="6397" lane="2" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Danuta" gender="F" lastname="Radkowiak" nation="POL" athleteid="1956">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="1957" heatid="6429" lane="4" entrytime="00:08:00.00" />
                <RESULT eventid="1183" points="406" reactiontime="+110" swimtime="00:04:00.88" resultid="1958" heatid="6105" lane="6" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.24" />
                    <SPLIT distance="100" swimtime="00:02:00.25" />
                    <SPLIT distance="150" swimtime="00:03:01.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="302" reactiontime="+106" swimtime="00:04:15.76" resultid="1959" heatid="6181" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.58" />
                    <SPLIT distance="100" swimtime="00:02:02.31" />
                    <SPLIT distance="150" swimtime="00:03:08.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" status="DNS" swimtime="00:00:00.00" resultid="1960" heatid="6294" lane="5" entrytime="00:03:50.00" />
                <RESULT eventid="1483" points="286" reactiontime="+103" swimtime="00:01:51.51" resultid="1961" heatid="6312" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="1962" heatid="6506" lane="4" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Barbara" gender="F" lastname="Chomicka" nation="POL" athleteid="1963">
              <RESULTS>
                <RESULT eventid="1058" points="344" reactiontime="+110" swimtime="00:09:07.73" resultid="1964" heatid="6429" lane="5" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.98" />
                    <SPLIT distance="100" swimtime="00:02:14.81" />
                    <SPLIT distance="150" swimtime="00:03:23.43" />
                    <SPLIT distance="200" swimtime="00:04:33.06" />
                    <SPLIT distance="250" swimtime="00:05:45.08" />
                    <SPLIT distance="300" swimtime="00:06:59.37" />
                    <SPLIT distance="350" swimtime="00:08:05.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="359" reactiontime="+110" swimtime="00:01:55.34" resultid="1965" heatid="6075" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="339" reactiontime="+114" swimtime="00:04:44.45" resultid="1966" heatid="6181" lane="4" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.69" />
                    <SPLIT distance="100" swimtime="00:02:17.42" />
                    <SPLIT distance="150" swimtime="00:03:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="253" reactiontime="+102" swimtime="00:00:57.85" resultid="1967" heatid="6219" lane="6" entrytime="00:00:55.00" />
                <RESULT eventid="1452" points="296" reactiontime="+110" swimtime="00:04:30.39" resultid="1968" heatid="6293" lane="3" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.94" />
                    <SPLIT distance="100" swimtime="00:02:13.15" />
                    <SPLIT distance="150" swimtime="00:03:25.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="249" reactiontime="+104" swimtime="00:02:10.96" resultid="1969" heatid="6312" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="350" reactiontime="+108" swimtime="00:02:02.57" resultid="1970" heatid="6505" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Hanka" gender="F" lastname="Kania" nation="POL" athleteid="1971">
              <RESULTS>
                <RESULT eventid="1153" points="441" reactiontime="+113" swimtime="00:01:41.76" resultid="1972" heatid="6076" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="556" reactiontime="+115" swimtime="00:03:50.87" resultid="1973" heatid="6104" lane="4" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.40" />
                    <SPLIT distance="100" swimtime="00:01:51.11" />
                    <SPLIT distance="150" swimtime="00:02:51.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="349" reactiontime="+111" swimtime="00:00:47.64" resultid="1974" heatid="6219" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="1422" points="437" reactiontime="+115" swimtime="00:03:18.23" resultid="1975" heatid="6274" lane="6" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:01:32.95" />
                    <SPLIT distance="150" swimtime="00:02:25.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="317" reactiontime="+115" swimtime="00:01:53.02" resultid="1976" heatid="6313" lane="5" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="451" reactiontime="+110" swimtime="00:01:53.77" resultid="1977" heatid="6507" lane="6" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1923-01-01" firstname="Danuta" gender="F" lastname="Kowalewska" nation="POL" athleteid="1978">
              <RESULTS>
                <RESULT eventid="1318" points="130" swimtime="00:02:15.85" resultid="1979" heatid="6192" lane="2" entrytime="00:01:48.00" />
                <RESULT eventid="1595" points="153" swimtime="00:05:04.33" resultid="1980" heatid="6503" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:40.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="1981">
              <RESULTS>
                <RESULT eventid="1198" points="542" reactiontime="+99" swimtime="00:03:58.96" resultid="1982" heatid="6110" lane="5" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.33" />
                    <SPLIT distance="100" swimtime="00:01:53.31" />
                    <SPLIT distance="150" swimtime="00:02:57.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="622" reactiontime="+99" swimtime="00:00:44.78" resultid="1983" heatid="6208" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1467" points="523" reactiontime="+104" swimtime="00:03:50.50" resultid="1984" heatid="6301" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.22" />
                    <SPLIT distance="100" swimtime="00:01:50.95" />
                    <SPLIT distance="150" swimtime="00:02:55.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="448" reactiontime="+104" swimtime="00:00:39.38" resultid="1985" heatid="6344" lane="2" entrytime="00:00:36.50" />
                <RESULT eventid="1610" points="553" reactiontime="+104" swimtime="00:01:46.60" resultid="1986" heatid="6397" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Renata" gender="F" lastname="Polańczyk" nation="POL" athleteid="1987">
              <RESULTS>
                <RESULT eventid="1058" points="374" reactiontime="+104" swimtime="00:08:05.46" resultid="1988" heatid="6429" lane="2" entrytime="00:08:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.31" />
                    <SPLIT distance="100" swimtime="00:01:53.20" />
                    <SPLIT distance="150" swimtime="00:02:48.16" />
                    <SPLIT distance="200" swimtime="00:03:43.13" />
                    <SPLIT distance="250" swimtime="00:05:00.49" />
                    <SPLIT distance="300" swimtime="00:06:19.04" />
                    <SPLIT distance="350" swimtime="00:07:15.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="346" reactiontime="+108" swimtime="00:01:47.66" resultid="1989" heatid="6076" lane="3" entrytime="00:01:44.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="377" reactiontime="+113" swimtime="00:03:57.39" resultid="1990" heatid="6182" lane="6" entrytime="00:03:59.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.95" />
                    <SPLIT distance="100" swimtime="00:01:55.05" />
                    <SPLIT distance="150" swimtime="00:02:57.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="512" reactiontime="+74" swimtime="00:01:36.49" resultid="1991" heatid="6245" lane="3" entrytime="00:01:35.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" status="DNS" swimtime="00:00:00.00" resultid="1992" heatid="6294" lane="2" entrytime="00:03:44.89" />
                <RESULT eventid="1543" points="517" reactiontime="+71" swimtime="00:03:33.18" resultid="1993" heatid="6369" lane="6" entrytime="00:03:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.38" />
                    <SPLIT distance="100" swimtime="00:01:45.60" />
                    <SPLIT distance="150" swimtime="00:02:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="435" reactiontime="+118" swimtime="00:06:47.74" resultid="1994" heatid="6555" lane="4" entrytime="00:06:42.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                    <SPLIT distance="100" swimtime="00:01:35.39" />
                    <SPLIT distance="150" swimtime="00:02:27.21" />
                    <SPLIT distance="200" swimtime="00:03:19.69" />
                    <SPLIT distance="250" swimtime="00:04:13.18" />
                    <SPLIT distance="300" swimtime="00:05:07.36" />
                    <SPLIT distance="350" swimtime="00:06:00.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Piotr" gender="M" lastname="Stasiuk" nation="POL" athleteid="1995">
              <RESULTS>
                <RESULT eventid="1168" points="472" reactiontime="+84" swimtime="00:01:19.24" resultid="1996" heatid="6092" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="561" reactiontime="+81" swimtime="00:00:32.31" resultid="1997" heatid="6233" lane="1" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Katarzyna" gender="F" lastname="Mazurek" nation="POL" athleteid="1998">
              <RESULTS>
                <RESULT eventid="1153" points="577" reactiontime="+110" swimtime="00:01:30.78" resultid="1999" heatid="6079" lane="6" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="495" reactiontime="+95" swimtime="00:01:22.18" resultid="2000" heatid="6153" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="701" swimtime="00:00:42.66" resultid="2001" heatid="6199" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1348" points="549" reactiontime="+92" swimtime="00:00:40.26" resultid="2002" heatid="6220" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1483" points="427" reactiontime="+91" swimtime="00:01:37.58" resultid="2003" heatid="6314" lane="2" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="501" reactiontime="+95" swimtime="00:00:36.68" resultid="2004" heatid="6336" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT comment="O-4 - przedwczesny start." eventid="1243" reactiontime="+71" status="DSQ" swimtime="00:02:50.85" resultid="1723" heatid="6519" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.30" />
                    <SPLIT distance="100" swimtime="00:01:28.58" />
                    <SPLIT distance="150" swimtime="00:02:14.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1987" number="1" reactiontime="+71" status="DSQ" />
                    <RELAYPOSITION athleteid="1943" number="2" reactiontime="+78" status="DSQ" />
                    <RELAYPOSITION athleteid="1998" number="3" reactiontime="+10" status="DSQ" />
                    <RELAYPOSITION athleteid="1956" number="4" reactiontime="-25" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1408" reactiontime="+104" swimtime="00:02:31.10" resultid="1724" heatid="6527" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                    <SPLIT distance="100" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:54.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1987" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="1943" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="1956" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="1998" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+76" swimtime="00:02:46.04" resultid="1722" heatid="6535" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                    <SPLIT distance="100" swimtime="00:01:29.83" />
                    <SPLIT distance="150" swimtime="00:02:10.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1987" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="1950" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="1998" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="1981" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1107" reactiontime="+110" swimtime="00:02:31.22" resultid="2005" heatid="6494" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                    <SPLIT distance="150" swimtime="00:01:53.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1950" number="1" reactiontime="+110" />
                    <RELAYPOSITION athleteid="1956" number="2" />
                    <RELAYPOSITION athleteid="1981" number="3" />
                    <RELAYPOSITION athleteid="1998" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Niezrzeszony Wrocław" nation="POL">
          <CONTACT name="asd" />
          <ATHLETES>
            <ATHLETE birthdate="1989-03-15" firstname="Bartłomiej" gender="M" lastname="Jankowski" nation="POL" athleteid="1731">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="1732" heatid="6490" lane="4" entrytime="00:06:04.00" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="1733" heatid="6117" lane="6" entrytime="00:02:40.00" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="1734" heatid="6188" lane="2" entrytime="00:03:00.00" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="1735" heatid="6215" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="1736" heatid="6306" lane="4" entrytime="00:02:49.00" />
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="1737" heatid="6379" lane="5" entrytime="00:02:43.00" />
                <RESULT eventid="1610" status="DNS" swimtime="00:00:00.00" resultid="1738" heatid="6406" lane="4" entrytime="00:01:16.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Niezrzeszony Jarosław" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Tomasz" gender="M" lastname="Jaroń" nation="POL" athleteid="1740">
              <RESULTS>
                <RESULT eventid="1092" points="427" reactiontime="+78" swimtime="00:06:29.60" resultid="1741" heatid="6489" lane="6" entrytime="00:06:21.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                    <SPLIT distance="100" swimtime="00:01:27.20" />
                    <SPLIT distance="150" swimtime="00:02:20.55" />
                    <SPLIT distance="200" swimtime="00:03:14.00" />
                    <SPLIT distance="250" swimtime="00:04:06.50" />
                    <SPLIT distance="300" swimtime="00:05:00.55" />
                    <SPLIT distance="350" swimtime="00:05:44.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="508" reactiontime="+79" swimtime="00:03:08.39" resultid="1742" heatid="6113" lane="5" entrytime="00:03:07.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.84" />
                    <SPLIT distance="100" swimtime="00:01:29.11" />
                    <SPLIT distance="150" swimtime="00:02:19.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="268" reactiontime="+79" swimtime="00:03:22.22" resultid="1743" heatid="6187" lane="3" entrytime="00:03:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:27.13" />
                    <SPLIT distance="150" swimtime="00:02:22.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="371" reactiontime="+77" swimtime="00:00:37.10" resultid="1744" heatid="6230" lane="6" entrytime="00:00:33.99" />
                <RESULT eventid="1467" points="424" reactiontime="+79" swimtime="00:03:01.41" resultid="1745" heatid="6304" lane="4" entrytime="00:02:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:27.43" />
                    <SPLIT distance="150" swimtime="00:02:19.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="1746" heatid="6351" lane="2" entrytime="00:00:30.99" />
                <RESULT eventid="1640" status="DNS" swimtime="00:00:00.00" resultid="1747" heatid="6565" lane="6" entrytime="00:05:36.99" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Konstancin-Jeziorna" nation="POL">
          <CONTACT name="Obiedziński" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-11" firstname="Paweł" gender="M" lastname="Obiedziński" nation="POL" athleteid="1749">
              <RESULTS>
                <RESULT eventid="1168" points="624" reactiontime="+78" swimtime="00:01:12.21" resultid="1750" heatid="6093" lane="3" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="671" reactiontime="+72" swimtime="00:01:01.01" resultid="1751" heatid="6173" lane="6" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="601" reactiontime="+75" swimtime="00:00:31.59" resultid="1752" heatid="6232" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="1437" points="626" reactiontime="+78" swimtime="00:02:18.34" resultid="1753" heatid="6288" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:06.40" />
                    <SPLIT distance="150" swimtime="00:01:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="708" reactiontime="+76" swimtime="00:00:27.39" resultid="1754" heatid="6356" lane="3" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="MKP Szczecin" nation="POL">
          <CONTACT city="Szczecin" email="windmuhle@wp.pl" name="Kowalczyk Piotr" phone="509758055" state="ZACH" street="Kaliny 45/9" zip="71-118" />
          <ATHLETES>
            <ATHLETE birthdate="1935-08-21" firstname="STEFANIA" gender="F" lastname="NOETZEL" nation="POL" athleteid="1757">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. K" eventid="1318" points="433" swimtime="00:01:02.31" resultid="6512" heatid="6192" lane="1" />
                <RESULT eventid="1595" points="568" swimtime="00:02:13.88" resultid="6513" heatid="6502" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.10" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="rekord Polski kat. K" eventid="1183" points="733" swimtime="00:04:42.66" resultid="6511" heatid="6101" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.49" />
                    <SPLIT distance="100" swimtime="00:02:21.25" />
                    <SPLIT distance="150" swimtime="00:03:33.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="2462">
              <RESULTS>
                <RESULT eventid="1137" points="589" swimtime="00:10:14.38" resultid="2463" heatid="6455" lane="5" entrytime="00:10:19.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="200" swimtime="00:02:25.12" />
                    <SPLIT distance="300" swimtime="00:03:42.62" />
                    <SPLIT distance="400" swimtime="00:05:00.66" />
                    <SPLIT distance="500" swimtime="00:06:18.91" />
                    <SPLIT distance="600" swimtime="00:07:38.82" />
                    <SPLIT distance="700" swimtime="00:08:58.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="626" reactiontime="+80" swimtime="00:01:00.11" resultid="2464" heatid="6174" lane="5" entrytime="00:01:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="659" reactiontime="+80" swimtime="00:02:13.45" resultid="2465" heatid="6289" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="100" swimtime="00:01:06.10" />
                    <SPLIT distance="150" swimtime="00:01:40.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="2466" heatid="6358" lane="5" entrytime="00:00:27.80" />
                <RESULT eventid="1640" points="622" reactiontime="+78" swimtime="00:04:47.50" resultid="2467" heatid="6567" lane="3" entrytime="00:04:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:08.63" />
                    <SPLIT distance="150" swimtime="00:01:44.82" />
                    <SPLIT distance="200" swimtime="00:02:22.15" />
                    <SPLIT distance="250" swimtime="00:02:59.12" />
                    <SPLIT distance="300" swimtime="00:03:36.20" />
                    <SPLIT distance="350" swimtime="00:04:12.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-08" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="2468">
              <RESULTS>
                <RESULT eventid="1257" points="854" reactiontime="+54" swimtime="00:01:06.96" resultid="2469" heatid="6157" lane="4" entrytime="00:01:07.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="870" swimtime="00:02:24.52" resultid="2470" heatid="6277" lane="2" entrytime="00:02:22.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:10.07" />
                    <SPLIT distance="150" swimtime="00:01:47.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="867" reactiontime="+73" swimtime="00:05:07.20" resultid="2471" heatid="6558" lane="3" entrytime="00:04:59.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:12.97" />
                    <SPLIT distance="150" swimtime="00:01:51.65" />
                    <SPLIT distance="200" swimtime="00:02:30.98" />
                    <SPLIT distance="250" swimtime="00:03:10.54" />
                    <SPLIT distance="300" swimtime="00:03:49.98" />
                    <SPLIT distance="350" swimtime="00:04:29.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="MOSiR  Częstochowa" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1969-01-01" firstname="Ireneusz" gender="M" lastname="Stachurski" nation="POL" athleteid="1762">
              <RESULTS>
                <RESULT eventid="1228" points="291" reactiontime="+82" swimtime="00:00:42.28" resultid="1763" heatid="6130" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1393" points="287" reactiontime="+79" swimtime="00:01:31.98" resultid="1764" heatid="6252" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="321" reactiontime="+74" swimtime="00:03:17.76" resultid="1765" heatid="6374" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                    <SPLIT distance="100" swimtime="00:01:34.76" />
                    <SPLIT distance="150" swimtime="00:02:26.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Niezrzeszeni" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1962-01-01" firstname="Mariola" gender="F" lastname="Strychalska" nation="POL" athleteid="1767">
              <RESULTS>
                <RESULT eventid="1213" points="471" reactiontime="+82" swimtime="00:00:44.47" resultid="1768" heatid="6121" lane="3" entrytime="00:00:44.93" />
                <RESULT eventid="1257" points="406" reactiontime="+113" swimtime="00:01:27.81" resultid="1769" heatid="6148" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="465" reactiontime="+113" swimtime="00:00:48.93" resultid="1770" heatid="6197" lane="1" entrytime="00:00:49.23" />
                <RESULT eventid="1378" points="509" reactiontime="+91" swimtime="00:01:36.68" resultid="1771" heatid="6242" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="438" reactiontime="+104" swimtime="00:00:38.35" resultid="1772" heatid="6333" lane="5" entrytime="00:00:38.37" />
                <RESULT eventid="1595" points="412" reactiontime="+114" swimtime="00:01:52.00" resultid="1773" heatid="6506" lane="3" entrytime="00:01:49.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Andrzej" gender="M" lastname="Chudy" nation="POL" athleteid="2063">
              <RESULTS>
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="2064" heatid="6449" lane="2" entrytime="00:13:20.76" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="2065" heatid="6133" lane="5" entrytime="00:00:35.94" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="2066" heatid="6160" lane="2" entrytime="00:01:32.99" />
                <RESULT eventid="1393" status="DNS" swimtime="00:00:00.00" resultid="2067" heatid="6253" lane="3" entrytime="00:01:31.75" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="2068" heatid="6285" lane="2" entrytime="00:02:31.23" />
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="2069" heatid="6375" lane="5" entrytime="00:03:22.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Arkadiusz" gender="M" lastname="Doliński" nation="POL" athleteid="2088">
              <RESULTS>
                <RESULT eventid="1228" points="510" reactiontime="+63" swimtime="00:00:32.66" resultid="2089" heatid="6135" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1393" points="445" reactiontime="+73" swimtime="00:01:14.20" resultid="2090" heatid="6258" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="2104">
              <RESULTS>
                <RESULT eventid="1228" points="575" reactiontime="+83" swimtime="00:00:38.37" resultid="2105" heatid="6131" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1272" points="540" reactiontime="+94" swimtime="00:01:12.03" resultid="2106" heatid="6164" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="445" reactiontime="+99" swimtime="00:01:28.49" resultid="2107" heatid="6254" lane="1" entrytime="00:01:30.00" />
                <RESULT eventid="1467" points="489" reactiontime="+95" swimtime="00:03:16.35" resultid="2108" heatid="6301" lane="2" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                    <SPLIT distance="100" swimtime="00:01:33.76" />
                    <SPLIT distance="150" swimtime="00:02:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="569" reactiontime="+88" swimtime="00:00:31.50" resultid="2109" heatid="6349" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1558" points="425" reactiontime="+88" swimtime="00:03:20.31" resultid="2110" heatid="6374" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.99" />
                    <SPLIT distance="150" swimtime="00:02:33.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1137" points="432" swimtime="00:13:14.84" resultid="6039" heatid="6448" lane="3" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:01:25.58" />
                    <SPLIT distance="200" swimtime="00:03:03.02" />
                    <SPLIT distance="300" swimtime="00:04:44.11" />
                    <SPLIT distance="400" swimtime="00:06:27.94" />
                    <SPLIT distance="500" swimtime="00:08:11.90" />
                    <SPLIT distance="600" swimtime="00:09:55.32" />
                    <SPLIT distance="700" swimtime="00:11:39.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Aleksandra" gender="F" lastname="Kącki" nation="POL" athleteid="2126">
              <RESULTS>
                <RESULT eventid="1513" points="287" reactiontime="+96" swimtime="00:00:41.22" resultid="2127" heatid="6331" lane="5" entrytime="00:00:43.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Wiesław" gender="M" lastname="Majcher" nation="POL" athleteid="2617">
              <RESULTS>
                <RESULT eventid="1137" points="183" swimtime="00:17:48.48" resultid="2618" heatid="6446" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.51" />
                    <SPLIT distance="100" swimtime="00:01:52.48" />
                    <SPLIT distance="200" swimtime="00:04:05.92" />
                    <SPLIT distance="300" swimtime="00:06:23.80" />
                    <SPLIT distance="400" swimtime="00:08:36.02" />
                    <SPLIT distance="500" swimtime="00:10:51.33" />
                    <SPLIT distance="600" swimtime="00:13:09.11" />
                    <SPLIT distance="700" swimtime="00:15:28.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="263" reactiontime="+88" swimtime="00:01:37.25" resultid="2619" heatid="6159" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="197" reactiontime="+116" swimtime="00:00:52.18" resultid="2620" heatid="6224" lane="1" />
                <RESULT eventid="1528" points="296" reactiontime="+61" swimtime="00:00:40.92" resultid="2621" heatid="6341" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1931-01-01" firstname="Jan" gender="M" lastname="Ślężyński" nation="POL" athleteid="2622">
              <RESULTS>
                <RESULT eventid="1137" points="258" swimtime="00:22:44.91" resultid="2623" heatid="6447" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.20" />
                    <SPLIT distance="100" swimtime="00:02:39.10" />
                    <SPLIT distance="200" swimtime="00:05:35.20" />
                    <SPLIT distance="300" swimtime="00:08:27.35" />
                    <SPLIT distance="400" swimtime="00:11:21.20" />
                    <SPLIT distance="500" swimtime="00:14:13.54" />
                    <SPLIT distance="600" swimtime="00:17:08.01" />
                    <SPLIT distance="700" swimtime="00:20:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="368" swimtime="00:05:39.72" resultid="2624" heatid="6108" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.37" />
                    <SPLIT distance="100" swimtime="00:02:43.21" />
                    <SPLIT distance="150" swimtime="00:04:11.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="218" swimtime="00:05:19.77" resultid="2625" heatid="6278" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.45" />
                    <SPLIT distance="100" swimtime="00:02:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="253" reactiontime="+74" swimtime="00:10:50.88" resultid="2626" heatid="6560" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.21" />
                    <SPLIT distance="100" swimtime="00:02:28.79" />
                    <SPLIT distance="150" swimtime="00:03:53.93" />
                    <SPLIT distance="200" swimtime="00:05:18.41" />
                    <SPLIT distance="250" swimtime="00:06:40.84" />
                    <SPLIT distance="300" swimtime="00:08:05.21" />
                    <SPLIT distance="350" swimtime="00:09:29.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-03" firstname="Konrad" gender="M" lastname="Gałka" nation="POL" athleteid="2847">
              <RESULTS>
                <RESULT eventid="1168" points="496" reactiontime="+92" swimtime="00:01:13.73" resultid="2848" heatid="6098" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="2849" heatid="6191" lane="6" entrytime="00:02:25.00" />
                <RESULT eventid="1363" points="567" reactiontime="+84" swimtime="00:00:30.36" resultid="2850" heatid="6239" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="2851" heatid="6310" lane="5" entrytime="00:02:30.00" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2852" heatid="6326" lane="2" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Anita" gender="F" lastname="Tworek" nation="POL" athleteid="2878">
              <RESULTS>
                <RESULT eventid="1122" points="204" swimtime="00:16:01.60" resultid="2879" heatid="6442" lane="6" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.34" />
                    <SPLIT distance="200" swimtime="00:03:50.06" />
                    <SPLIT distance="300" swimtime="00:05:53.64" />
                    <SPLIT distance="400" swimtime="00:07:52.96" />
                    <SPLIT distance="500" swimtime="00:09:55.28" />
                    <SPLIT distance="600" swimtime="00:11:57.70" />
                    <SPLIT distance="700" swimtime="00:14:01.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="137" reactiontime="+97" swimtime="00:01:00.94" resultid="2880" heatid="6120" lane="4" entrytime="00:00:54.00" />
                <RESULT eventid="1257" points="182" reactiontime="+102" swimtime="00:01:44.02" resultid="2881" heatid="6150" lane="1" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="188" reactiontime="+100" swimtime="00:00:59.38" resultid="2882" heatid="6194" lane="3" entrytime="00:00:54.00" />
                <RESULT eventid="1378" points="130" reactiontime="+87" swimtime="00:02:11.61" resultid="2883" heatid="6244" lane="4" entrytime="00:02:00.00" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="2884" heatid="6331" lane="1" entrytime="00:00:44.00" />
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="2885" heatid="6504" lane="3" entrytime="00:02:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Maria" gender="F" lastname="Ochab" nation="POL" athleteid="2886">
              <RESULTS>
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="2887" heatid="6120" lane="2" entrytime="00:00:54.00" />
                <RESULT eventid="1257" status="DNS" swimtime="00:00:00.00" resultid="2888" heatid="6150" lane="5" entrytime="00:01:42.00" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="2889" heatid="6195" lane="6" entrytime="00:00:54.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="2890" heatid="6272" lane="6" entrytime="00:03:46.00" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="2891" heatid="6331" lane="4" entrytime="00:00:43.00" />
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="2892" heatid="6505" lane="6" entrytime="00:02:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Piotr" gender="M" lastname="Kalinowski" nation="POL" athleteid="2893">
              <RESULTS>
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="2894" heatid="6454" lane="4" entrytime="00:10:33.70" />
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="2895" heatid="6095" lane="1" entrytime="00:01:10.98" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="2896" heatid="6173" lane="3" entrytime="00:01:00.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Hanna" gender="F" lastname="Rutkowska" nation="POL" athleteid="3288">
              <RESULTS>
                <RESULT eventid="1513" points="496" reactiontime="+87" swimtime="00:00:32.34" resultid="3289" heatid="6337" lane="3" entrytime="00:00:32.05" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Artur" gender="M" lastname="Wszołek" nation="POL" athleteid="3290">
              <RESULTS>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="3291" heatid="6170" lane="4" entrytime="00:01:05.00" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3292" heatid="6352" lane="3" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Krystyna" gender="F" lastname="Tokarska" nation="POL" athleteid="3293">
              <RESULTS>
                <RESULT eventid="1122" points="213" swimtime="00:15:47.77" resultid="3294" heatid="6441" lane="3" entrytime="00:16:15.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                    <SPLIT distance="100" swimtime="00:01:43.84" />
                    <SPLIT distance="200" swimtime="00:03:43.48" />
                    <SPLIT distance="300" swimtime="00:05:45.72" />
                    <SPLIT distance="400" swimtime="00:07:47.44" />
                    <SPLIT distance="500" swimtime="00:09:46.79" />
                    <SPLIT distance="600" swimtime="00:11:49.16" />
                    <SPLIT distance="700" swimtime="00:13:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="319" reactiontime="+112" swimtime="00:03:58.94" resultid="3295" heatid="6104" lane="1" entrytime="00:04:01.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.13" />
                    <SPLIT distance="100" swimtime="00:01:52.36" />
                    <SPLIT distance="150" swimtime="00:02:56.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="206" reactiontime="+70" swimtime="00:00:53.16" resultid="3296" heatid="6119" lane="3" entrytime="00:00:58.30" />
                <RESULT eventid="1378" points="161" reactiontime="+73" swimtime="00:02:02.36" resultid="3297" heatid="6244" lane="1" entrytime="00:02:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="222" reactiontime="+101" swimtime="00:03:34.30" resultid="3298" heatid="6272" lane="3" entrytime="00:03:37.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                    <SPLIT distance="100" swimtime="00:01:38.85" />
                    <SPLIT distance="150" swimtime="00:02:37.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="173" reactiontime="+75" swimtime="00:04:20.72" resultid="3299" heatid="6367" lane="4" entrytime="00:04:20.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.47" />
                    <SPLIT distance="100" swimtime="00:02:07.74" />
                    <SPLIT distance="150" swimtime="00:03:15.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="206" reactiontime="+110" swimtime="00:07:40.40" resultid="3300" heatid="6554" lane="3" entrytime="00:07:34.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                    <SPLIT distance="100" swimtime="00:01:43.68" />
                    <SPLIT distance="150" swimtime="00:02:43.18" />
                    <SPLIT distance="200" swimtime="00:03:43.84" />
                    <SPLIT distance="250" swimtime="00:04:43.48" />
                    <SPLIT distance="300" swimtime="00:05:42.57" />
                    <SPLIT distance="350" swimtime="00:06:42.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Anna" gender="F" lastname="Spieszny" nation="POL" athleteid="3520">
              <RESULTS>
                <RESULT eventid="1318" points="291" reactiontime="+105" swimtime="00:00:54.42" resultid="3521" heatid="6195" lane="1" entrytime="00:00:53.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-11-21" firstname="Zbigniew" gender="M" lastname="Dymecki" nation="POL" athleteid="3851">
              <RESULTS>
                <RESULT eventid="1092" points="344" reactiontime="+110" swimtime="00:09:24.80" resultid="3852" heatid="6485" lane="1" entrytime="00:09:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.47" />
                    <SPLIT distance="100" swimtime="00:02:21.95" />
                    <SPLIT distance="150" swimtime="00:03:39.15" />
                    <SPLIT distance="200" swimtime="00:04:50.91" />
                    <SPLIT distance="250" swimtime="00:06:05.93" />
                    <SPLIT distance="300" swimtime="00:07:20.09" />
                    <SPLIT distance="350" swimtime="00:08:22.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="273" reactiontime="+105" swimtime="00:01:58.91" resultid="3853" heatid="6084" lane="6" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="236" reactiontime="+104" swimtime="00:05:12.83" resultid="3854" heatid="6183" lane="2" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.47" />
                    <SPLIT distance="100" swimtime="00:02:27.02" />
                    <SPLIT distance="150" swimtime="00:03:49.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="307" swimtime="00:00:50.56" resultid="3855" heatid="6224" lane="2" entrytime="00:00:52.00" />
                <RESULT eventid="1467" points="415" reactiontime="+112" swimtime="00:04:08.96" resultid="3856" heatid="6300" lane="1" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                    <SPLIT distance="100" swimtime="00:01:57.87" />
                    <SPLIT distance="150" swimtime="00:03:08.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="246" reactiontime="+125" swimtime="00:02:08.47" resultid="3857" heatid="6316" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="284" reactiontime="+108" swimtime="00:08:27.89" resultid="3858" heatid="6560" lane="4" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.69" />
                    <SPLIT distance="150" swimtime="00:02:53.33" />
                    <SPLIT distance="200" swimtime="00:04:00.99" />
                    <SPLIT distance="250" swimtime="00:05:09.54" />
                    <SPLIT distance="300" swimtime="00:06:17.44" />
                    <SPLIT distance="350" swimtime="00:07:22.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Jarosław" gender="M" lastname="Wyrwa" nation="POL" athleteid="3883">
              <RESULTS>
                <RESULT comment="O-4 - przedwczesny start." eventid="1333" reactiontime="+57" status="DSQ" swimtime="00:00:38.26" resultid="3884" heatid="6211" lane="3" entrytime="00:00:37.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Tomasz" gender="M" lastname="Stefaniak" nation="POL" athleteid="3885">
              <RESULTS>
                <RESULT eventid="1363" status="DNS" swimtime="00:00:00.00" resultid="3886" heatid="6230" lane="3" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Przemysław" gender="M" lastname="Kuśmider" nation="POL" athleteid="3887">
              <RESULTS>
                <RESULT eventid="1437" points="296" reactiontime="+86" swimtime="00:02:41.48" resultid="3888" heatid="6291" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:13.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Tomasz" gender="M" lastname="Zembala" nation="POL" athleteid="3889">
              <RESULTS>
                <RESULT comment="Z2" eventid="1168" reactiontime="+106" status="DSQ" swimtime="00:01:24.20" resultid="3891" heatid="6087" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="417" reactiontime="+100" swimtime="00:01:11.46" resultid="3892" heatid="6166" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="361" reactiontime="+103" swimtime="00:00:37.42" resultid="3893" heatid="6229" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="3894" heatid="6302" lane="2" entrytime="00:03:30.00" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="3895" heatid="6318" lane="5" entrytime="00:01:35.00" />
                <RESULT eventid="1528" points="453" reactiontime="+97" swimtime="00:00:31.79" resultid="3896" heatid="6351" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1137" points="386" swimtime="00:11:50.44" resultid="6038" heatid="6452" lane="6" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:19.81" />
                    <SPLIT distance="200" swimtime="00:02:48.97" />
                    <SPLIT distance="300" swimtime="00:04:18.66" />
                    <SPLIT distance="400" swimtime="00:05:50.53" />
                    <SPLIT distance="500" swimtime="00:07:22.34" />
                    <SPLIT distance="600" swimtime="00:08:53.59" />
                    <SPLIT distance="700" swimtime="00:10:23.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-06-07" firstname="Olga" gender="F" lastname="Krysiak" nation="POL" athleteid="3923">
              <RESULTS>
                <RESULT eventid="1257" points="666" reactiontime="+79" swimtime="00:01:03.91" resultid="3924" heatid="6158" lane="4" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="650" reactiontime="+78" swimtime="00:02:23.15" resultid="3925" heatid="6277" lane="5" entrytime="00:02:23.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:08.84" />
                    <SPLIT distance="150" swimtime="00:01:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="615" reactiontime="+78" swimtime="00:00:30.11" resultid="3926" heatid="6339" lane="3" entrytime="00:00:29.95" entrycourse="SCM" />
                <RESULT eventid="1625" points="525" reactiontime="+80" swimtime="00:05:14.31" resultid="3927" heatid="6558" lane="1" entrytime="00:05:12.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:12.91" />
                    <SPLIT distance="150" swimtime="00:01:52.78" />
                    <SPLIT distance="200" swimtime="00:02:32.79" />
                    <SPLIT distance="250" swimtime="00:03:13.38" />
                    <SPLIT distance="300" swimtime="00:03:54.23" />
                    <SPLIT distance="350" swimtime="00:04:35.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-17" firstname="Artur" gender="M" lastname="Włoszek" nation="POL" athleteid="4765">
              <RESULTS>
                <RESULT eventid="1272" points="587" reactiontime="+71" swimtime="00:01:00.49" resultid="4766" heatid="6167" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="651" reactiontime="+71" swimtime="00:00:26.61" resultid="4767" heatid="6353" lane="1" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-21" firstname="Ewelina " gender="F" lastname="Kot" nation="POL" athleteid="6028">
              <RESULTS>
                <RESULT eventid="1122" points="457" swimtime="00:11:20.86" resultid="6029" heatid="6445" lane="5" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:20.97" />
                    <SPLIT distance="150" swimtime="00:02:46.31" />
                    <SPLIT distance="200" swimtime="00:04:12.48" />
                    <SPLIT distance="300" swimtime="00:04:12.48" />
                    <SPLIT distance="400" swimtime="00:05:38.81" />
                    <SPLIT distance="500" swimtime="00:07:04.49" />
                    <SPLIT distance="600" swimtime="00:08:30.08" />
                    <SPLIT distance="700" swimtime="00:09:56.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Tarnowskie WOPR" nation="POL" region="MAL">
          <CONTACT city="zgłobice" name="kacer" phone="607681313" street="rzemieślnicza 24" zip="33-113" />
          <ATHLETES>
            <ATHLETE birthdate="1976-06-18" firstname="Paweł" gender="M" lastname="Pastuszko" nation="POL" athleteid="1775">
              <RESULTS>
                <RESULT eventid="1272" points="177" reactiontime="+95" swimtime="00:01:31.46" resultid="1776" heatid="6161" lane="5" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="150" reactiontime="+106" swimtime="00:03:38.56" resultid="1777" heatid="6282" lane="4" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:01:37.49" />
                    <SPLIT distance="150" swimtime="00:02:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="208" reactiontime="+104" swimtime="00:00:39.03" resultid="1778" heatid="6345" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-11" firstname="Przemysław" gender="M" lastname="Jurek" nation="POL" athleteid="1779">
              <RESULTS>
                <RESULT eventid="1137" status="DNF" swimtime="00:00:00.00" resultid="1780" heatid="6456" lane="4" entrytime="00:09:50.00" />
                <RESULT eventid="1168" points="579" reactiontime="+76" swimtime="00:01:09.89" resultid="1781" heatid="6098" lane="3" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="541" reactiontime="+80" swimtime="00:02:16.98" resultid="1782" heatid="6292" lane="1" entrytime="00:02:04.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                    <SPLIT distance="100" swimtime="00:01:03.69" />
                    <SPLIT distance="150" swimtime="00:01:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="479" reactiontime="+83" swimtime="00:05:07.41" resultid="1783" heatid="6570" lane="6" entrytime="00:04:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:09.43" />
                    <SPLIT distance="150" swimtime="00:01:48.93" />
                    <SPLIT distance="200" swimtime="00:02:28.76" />
                    <SPLIT distance="250" swimtime="00:03:09.16" />
                    <SPLIT distance="300" swimtime="00:03:49.14" />
                    <SPLIT distance="350" swimtime="00:04:29.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-15" firstname="Marcin" gender="M" lastname="Kacer" nation="POL" athleteid="1784">
              <RESULTS>
                <RESULT eventid="1272" points="595" reactiontime="+82" swimtime="00:01:00.21" resultid="1785" heatid="6179" lane="1" entrytime="00:00:56.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="712" reactiontime="+81" swimtime="00:00:28.28" resultid="1786" heatid="6241" lane="5" entrytime="00:00:26.99" />
                <RESULT eventid="1498" points="685" reactiontime="+82" swimtime="00:01:03.19" resultid="1787" heatid="6326" lane="4" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01711" name="UKS WODNIK Siemianowice Śląskie" nation="POL" region="SLA" shortname="UKS WODNIK Siemianowice Śląski">
          <CONTACT city="Siemianowice Śląskie" email="vivisektor@interia.pl" name="Małyszek Leszek" phone="534039934" state="SLA" street="Mikołaja 3" zip="41-106" />
          <ATHLETES>
            <ATHLETE birthdate="1981-06-06" firstname="Leszek" gender="M" lastname="Małyszek" nation="POL" athleteid="1789">
              <RESULTS>
                <RESULT eventid="1333" points="609" reactiontime="+59" swimtime="00:00:34.74" resultid="1790" heatid="6214" lane="2" entrytime="00:00:34.50" />
                <RESULT eventid="1610" points="554" reactiontime="+83" swimtime="00:01:18.95" resultid="1791" heatid="6405" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-08-05" firstname="Mateusz" gender="M" lastname="Miodoński" nation="POL" athleteid="1792">
              <RESULTS>
                <RESULT eventid="1168" points="582" reactiontime="+77" swimtime="00:01:09.33" resultid="1793" heatid="6099" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-07-28" firstname="Wojciech" gender="M" lastname="Zych" nation="POL" athleteid="1794">
              <RESULTS>
                <RESULT eventid="1333" points="709" reactiontime="+92" swimtime="00:00:37.23" resultid="1795" heatid="6213" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1363" points="676" reactiontime="+97" swimtime="00:00:31.98" resultid="1796" heatid="6234" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1528" points="638" reactiontime="+95" swimtime="00:00:30.33" resultid="1797" heatid="6352" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1610" status="DNS" swimtime="00:00:00.00" resultid="1798" heatid="6403" lane="2" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="1799">
              <RESULTS>
                <RESULT eventid="1137" points="567" swimtime="00:11:24.98" resultid="1800" heatid="6453" lane="5" entrytime="00:11:20.44">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.80" />
                    <SPLIT distance="200" swimtime="00:02:46.45" />
                    <SPLIT distance="300" swimtime="00:04:13.09" />
                    <SPLIT distance="400" swimtime="00:05:38.69" />
                    <SPLIT distance="500" swimtime="00:07:05.26" />
                    <SPLIT distance="600" swimtime="00:08:32.09" />
                    <SPLIT distance="700" swimtime="00:09:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="1801" heatid="6091" lane="4" entrytime="00:01:18.12" />
                <RESULT eventid="1302" points="424" reactiontime="+85" swimtime="00:03:19.89" resultid="1802" heatid="6187" lane="1" entrytime="00:03:11.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.94" />
                    <SPLIT distance="100" swimtime="00:01:33.55" />
                    <SPLIT distance="150" swimtime="00:02:26.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="488" reactiontime="+81" swimtime="00:00:35.22" resultid="1803" heatid="6228" lane="3" entrytime="00:00:35.20" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="1804" heatid="6305" lane="2" entrytime="00:02:52.30" />
                <RESULT eventid="1498" points="430" reactiontime="+81" swimtime="00:01:23.67" resultid="1805" heatid="6320" lane="4" entrytime="00:01:20.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="458" reactiontime="+81" swimtime="00:05:48.01" resultid="1806" heatid="6565" lane="3" entrytime="00:05:28.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                    <SPLIT distance="150" swimtime="00:02:06.03" />
                    <SPLIT distance="200" swimtime="00:02:50.66" />
                    <SPLIT distance="250" swimtime="00:03:35.45" />
                    <SPLIT distance="300" swimtime="00:04:20.69" />
                    <SPLIT distance="350" swimtime="00:05:05.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+63" swimtime="00:02:12.21" resultid="1807" heatid="6525" lane="1" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:06.72" />
                    <SPLIT distance="150" swimtime="00:01:42.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1792" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="1789" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="1799" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="1794" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Masters Płońsk" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1940-01-01" firstname="Wieczorkiewicz" gender="F" lastname="Alina" nation="POL" athleteid="1812">
              <RESULTS>
                <RESULT eventid="1153" points="158" reactiontime="+144" swimtime="00:02:58.52" resultid="1813" heatid="6074" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="175" reactiontime="+80" swimtime="00:01:17.82" resultid="1814" heatid="6118" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1318" points="130" reactiontime="+113" swimtime="00:01:27.72" resultid="1815" heatid="6192" lane="4" entrytime="00:01:45.00" />
                <RESULT comment="O4 - przedwczesny start," eventid="1378" reactiontime="+51" status="DSQ" swimtime="00:02:57.18" resultid="1816" heatid="6243" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="190" reactiontime="+88" swimtime="00:06:20.42" resultid="1817" heatid="6366" lane="3" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.98" />
                    <SPLIT distance="100" swimtime="00:03:04.67" />
                    <SPLIT distance="150" swimtime="00:04:52.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="148" reactiontime="+124" swimtime="00:03:08.56" resultid="1818" heatid="6503" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:32.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01805" name="Z-Ł Wopr Ozorków" nation="POL" region="LOD">
          <CONTACT city="OZORKÓW" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="LOTNICZA 1 A" zip="95-035" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-13" firstname="MIROSŁAWA" gender="F" lastname="RAJTAR" nation="POL" license="M0180510004" athleteid="1820">
              <RESULTS>
                <RESULT eventid="1153" points="541" reactiontime="+95" swimtime="00:01:35.06" resultid="1821" heatid="6078" lane="6" entrytime="00:01:37.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="507" reactiontime="+97" swimtime="00:01:25.92" resultid="1822" heatid="6152" lane="3" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="470" swimtime="00:00:43.14" resultid="1823" heatid="6219" lane="2" entrytime="00:00:47.40" entrycourse="SCM" />
                <RESULT eventid="1422" points="469" reactiontime="+89" swimtime="00:03:13.62" resultid="1824" heatid="6274" lane="1" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                    <SPLIT distance="100" swimtime="00:01:29.59" />
                    <SPLIT distance="150" swimtime="00:02:21.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="568" reactiontime="+96" swimtime="00:00:37.44" resultid="1825" heatid="6333" lane="4" entrytime="00:00:37.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="ROMAN" gender="M" lastname="WICZEL" nation="POL" license="M0180520003" athleteid="1826">
              <RESULTS>
                <RESULT eventid="1198" points="646" reactiontime="+98" swimtime="00:03:24.12" resultid="1827" heatid="6111" lane="2" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                    <SPLIT distance="100" swimtime="00:01:39.50" />
                    <SPLIT distance="150" swimtime="00:02:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="602" reactiontime="+86" swimtime="00:00:40.56" resultid="1828" heatid="6209" lane="4" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1610" points="697" reactiontime="+90" swimtime="00:01:29.09" resultid="1829" heatid="6400" lane="4" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-20" firstname="BOGDAN" gender="M" lastname="WĄSIK" nation="POL" license="M0180520002" athleteid="1830">
              <RESULTS>
                <RESULT eventid="1198" points="662" reactiontime="+93" swimtime="00:03:08.99" resultid="1831" heatid="6112" lane="3" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:01:29.75" />
                    <SPLIT distance="150" swimtime="00:02:19.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="1832" heatid="6186" lane="1" entrytime="00:03:34.00" entrycourse="SCM" />
                <RESULT eventid="1333" points="551" reactiontime="+96" swimtime="00:00:40.49" resultid="1833" heatid="6211" lane="6" entrytime="00:00:39.00" entrycourse="SCM" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="1834" heatid="6303" lane="5" entrytime="00:03:15.00" entrycourse="SCM" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="1835" heatid="6318" lane="2" entrytime="00:01:33.00" entrycourse="SCM" />
                <RESULT eventid="1610" points="617" reactiontime="+90" swimtime="00:01:27.25" resultid="1836" heatid="6402" lane="1" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="URSZULA" gender="F" lastname="MRÓZ" nation="POL" license="M0180510002" athleteid="1837">
              <RESULTS>
                <RESULT eventid="1153" points="695" reactiontime="+95" swimtime="00:01:25.33" resultid="1838" heatid="6079" lane="3" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. F" eventid="1213" points="736" reactiontime="+68" swimtime="00:00:38.32" resultid="1839" heatid="6124" lane="6" entrytime="00:00:38.50" entrycourse="SCM" />
                <RESULT eventid="1348" points="695" reactiontime="+99" swimtime="00:00:37.23" resultid="1840" heatid="6221" lane="5" entrytime="00:00:36.40" entrycourse="SCM" />
                <RESULT eventid="1513" points="653" reactiontime="+95" swimtime="00:00:33.58" resultid="1841" heatid="6336" lane="4" entrytime="00:00:33.70" entrycourse="SCM" />
                <RESULT eventid="1543" points="712" reactiontime="+65" swimtime="00:03:11.57" resultid="1842" heatid="6369" lane="4" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:28.26" />
                    <SPLIT distance="150" swimtime="00:02:19.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="EWA" gender="F" lastname="STĘPIEŃ" nation="POL" license="M0180510003" athleteid="1843">
              <RESULTS>
                <RESULT eventid="1153" points="699" reactiontime="+83" swimtime="00:01:25.19" resultid="1844" heatid="6080" lane="6" entrytime="00:01:24.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="635" reactiontime="+82" swimtime="00:01:15.64" resultid="1845" heatid="6154" lane="4" entrytime="00:01:15.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="801" reactiontime="+70" swimtime="00:00:40.82" resultid="1846" heatid="6200" lane="6" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1513" points="689" reactiontime="+73" swimtime="00:00:32.99" resultid="1847" heatid="6337" lane="6" entrytime="00:00:33.50" entrycourse="SCM" />
                <RESULT eventid="1595" points="769" reactiontime="+72" swimtime="00:01:30.96" resultid="1848" heatid="6509" lane="4" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="ZBIGNIEW" gender="M" lastname="MACIEJCZYK" nation="POL" license="M01805200" athleteid="1849">
              <RESULTS>
                <RESULT eventid="1272" points="654" reactiontime="+99" swimtime="00:01:16.07" resultid="1850" heatid="6162" lane="4" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="397" reactiontime="+102" swimtime="00:04:09.70" resultid="1851" heatid="6185" lane="4" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.04" />
                    <SPLIT distance="100" swimtime="00:01:55.76" />
                    <SPLIT distance="150" swimtime="00:03:05.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="575" reactiontime="+98" swimtime="00:00:38.30" resultid="1852" heatid="6228" lane="1" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1498" points="397" reactiontime="+103" swimtime="00:01:43.46" resultid="1853" heatid="6318" lane="4" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="638" reactiontime="+101" swimtime="00:00:32.83" resultid="1854" heatid="6344" lane="3" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-02-07" firstname="KRZYSZTOF" gender="M" lastname="WOJCIECHOWSKI" nation="POL" license="M01805200" athleteid="1855" />
            <ATHLETE birthdate="1957-01-09" firstname="WŁODZIMIERZ" gender="M" lastname="PRZYTULSKI" nation="POL" license="M0180520005" athleteid="1856">
              <RESULTS>
                <RESULT eventid="1228" points="712" reactiontime="+75" swimtime="00:00:35.72" resultid="1857" heatid="6133" lane="4" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1302" points="501" reactiontime="+89" swimtime="00:03:11.60" resultid="1858" heatid="6189" lane="6" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:28.00" />
                    <SPLIT distance="150" swimtime="00:02:20.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="637" reactiontime="+92" swimtime="00:00:32.62" resultid="1859" heatid="6232" lane="1" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="1860" heatid="6305" lane="4" entrytime="00:02:52.00" entrycourse="SCM" />
                <RESULT eventid="1498" points="519" reactiontime="+90" swimtime="00:01:20.05" resultid="1861" heatid="6321" lane="4" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1922-01-04" firstname="KAZIMIERZ" gender="M" lastname="MRÓWCZYŃSKI" nation="POL" license="M01805200" athleteid="1862">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. N" eventid="1137" points="883" swimtime="00:21:30.46" resultid="1863" heatid="6447" lane="5" entrytime="00:21:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:26.60" />
                    <SPLIT distance="200" swimtime="00:05:09.88" />
                    <SPLIT distance="300" swimtime="00:07:51.22" />
                    <SPLIT distance="400" swimtime="00:10:33.41" />
                    <SPLIT distance="500" swimtime="00:13:16.07" />
                    <SPLIT distance="600" swimtime="00:16:00.02" />
                    <SPLIT distance="700" swimtime="00:18:45.14" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. N" eventid="1272" points="654" reactiontime="+124" swimtime="00:02:08.25" resultid="1864" heatid="6159" lane="4" entrytime="00:02:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.94" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. N" eventid="1437" points="865" swimtime="00:04:46.07" resultid="1865" heatid="6278" lane="2" entrytime="00:04:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.09" />
                    <SPLIT distance="100" swimtime="00:02:17.26" />
                    <SPLIT distance="150" swimtime="00:03:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. N" eventid="1528" points="567" reactiontime="+121" swimtime="00:00:53.70" resultid="1866" heatid="6342" lane="2" entrytime="00:00:51.50" entrycourse="SCM" />
                <RESULT comment="Rekord Polski kat. N" eventid="1640" status="DNS" swimtime="00:00:00.00" resultid="1867" heatid="6560" lane="2" entrytime="00:10:20.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-07-18" firstname="TOMASZ" gender="M" lastname="NIEDZWIEDZ" nation="POL" license="M01805200" athleteid="1868">
              <RESULTS>
                <RESULT eventid="1092" points="361" reactiontime="+95" swimtime="00:07:06.29" resultid="1869" heatid="6487" lane="2" entrytime="00:07:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                    <SPLIT distance="100" swimtime="00:01:40.69" />
                    <SPLIT distance="150" swimtime="00:02:39.84" />
                    <SPLIT distance="200" swimtime="00:03:34.86" />
                    <SPLIT distance="250" swimtime="00:04:33.17" />
                    <SPLIT distance="300" swimtime="00:05:30.97" />
                    <SPLIT distance="350" swimtime="00:06:19.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="281" reactiontime="+62" swimtime="00:03:36.45" resultid="1870" heatid="6185" lane="2" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.27" />
                    <SPLIT distance="100" swimtime="00:01:42.04" />
                    <SPLIT distance="150" swimtime="00:02:39.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="1871" heatid="6302" lane="3" entrytime="00:03:25.00" entrycourse="SCM" />
                <RESULT eventid="1498" points="235" reactiontime="+103" swimtime="00:01:39.33" resultid="1872" heatid="6318" lane="6" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="340" reactiontime="+111" swimtime="00:01:38.47" resultid="1873" heatid="6397" lane="6" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-08" firstname="EWA" gender="F" lastname="ZIMNA-WALENDZIK" nation="POL" license="M0180510005" athleteid="1874">
              <RESULTS>
                <RESULT eventid="1153" points="530" reactiontime="+96" swimtime="00:01:41.32" resultid="1875" heatid="6076" lane="4" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="483" reactiontime="+89" swimtime="00:01:30.97" resultid="1876" heatid="6151" lane="5" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="438" reactiontime="+87" swimtime="00:00:48.17" resultid="1877" heatid="6219" lane="3" entrytime="00:00:45.00" entrycourse="SCM" />
                <RESULT eventid="1483" points="386" reactiontime="+89" swimtime="00:01:53.22" resultid="1878" heatid="6313" lane="1" entrytime="00:01:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="448" reactiontime="+86" swimtime="00:00:42.01" resultid="1879" heatid="6333" lane="6" entrytime="00:00:39.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-23" firstname="TOMASZ" gender="M" lastname="CAJDLER" nation="POL" license="M0180520006" athleteid="1880">
              <RESULTS>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="1881" heatid="6111" lane="1" entrytime="00:03:40.00" entrycourse="SCM" />
                <RESULT eventid="1272" points="509" reactiontime="+86" swimtime="00:01:11.25" resultid="1882" heatid="6165" lane="3" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="459" swimtime="00:00:41.74" resultid="1883" heatid="6209" lane="2" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1528" points="532" reactiontime="+91" swimtime="00:00:31.31" resultid="1884" heatid="6348" lane="6" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1610" points="432" reactiontime="+94" swimtime="00:01:36.26" resultid="1885" heatid="6400" lane="5" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+79" swimtime="00:02:30.86" resultid="1891" heatid="6523" lane="1" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:19.47" />
                    <SPLIT distance="150" swimtime="00:01:59.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1856" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="1830" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="1868" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="1880" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1415" swimtime="00:02:14.22" resultid="1892" heatid="6531" lane="4" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:07.20" />
                    <SPLIT distance="150" swimtime="00:01:43.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1880" number="1" />
                    <RELAYPOSITION athleteid="1868" number="2" />
                    <RELAYPOSITION athleteid="1830" number="3" />
                    <RELAYPOSITION athleteid="1856" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="2">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. E" eventid="1250" reactiontime="+86" swimtime="00:02:59.84" resultid="1893" heatid="6522" lane="2" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                    <SPLIT distance="100" swimtime="00:01:23.94" />
                    <SPLIT distance="150" swimtime="00:02:03.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1855" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="1826" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="1849" number="3" reactiontime="+92" />
                    <RELAYPOSITION athleteid="1862" number="4" reactiontime="+82" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1415" reactiontime="+100" swimtime="00:02:44.04" resultid="1894" heatid="6530" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.32" />
                    <SPLIT distance="100" swimtime="00:01:41.12" />
                    <SPLIT distance="150" swimtime="00:02:10.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1862" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="1826" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="1855" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="1849" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1243" reactiontime="+65" swimtime="00:02:43.14" resultid="1886" heatid="6520" lane="6" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                    <SPLIT distance="100" swimtime="00:01:25.76" />
                    <SPLIT distance="150" swimtime="00:02:02.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1820" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="1843" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="1837" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="1874" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1408" reactiontime="+93" swimtime="00:02:25.72" resultid="1888" heatid="6527" lane="3" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:01:52.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1837" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="1874" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="1820" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="1843" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Przedwczesny start." eventid="1107" reactiontime="+90" status="DSQ" swimtime="00:02:22.75" resultid="1889" heatid="6495" lane="3" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.90" />
                    <SPLIT distance="100" swimtime="00:01:51.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1820" number="1" reactiontime="+90" status="DSQ" />
                    <RELAYPOSITION athleteid="1855" number="2" reactiontime="+45" status="DSQ" />
                    <RELAYPOSITION athleteid="1874" number="3" reactiontime="-7" status="DSQ" />
                    <RELAYPOSITION athleteid="1849" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+76" swimtime="00:02:24.73" resultid="1895" heatid="6537" lane="1" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                    <SPLIT distance="150" swimtime="00:01:51.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1837" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="1830" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="1856" number="3" reactiontime="+73" />
                    <RELAYPOSITION athleteid="1843" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+67" swimtime="00:02:45.85" resultid="1890" heatid="6536" lane="4" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.60" />
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                    <SPLIT distance="150" swimtime="00:02:05.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1820" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="1826" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="1849" number="3" reactiontime="+95" />
                    <RELAYPOSITION athleteid="1874" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+79" swimtime="00:02:08.11" resultid="1942" heatid="6496" lane="4" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="150" swimtime="00:01:35.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1856" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="1837" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="1880" number="3" />
                    <RELAYPOSITION athleteid="1843" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="WOPR Tczew" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1987-01-01" firstname="Hebel" gender="F" lastname="Aleksandra" nation="POL" athleteid="1920">
              <RESULTS>
                <RESULT eventid="1213" points="352" reactiontime="+88" swimtime="00:00:43.10" resultid="1921" heatid="6123" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="1257" points="431" reactiontime="+83" swimtime="00:01:16.06" resultid="1922" heatid="6155" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" status="DNS" swimtime="00:00:00.00" resultid="1923" heatid="6246" lane="4" entrytime="00:01:31.00" />
                <RESULT eventid="1422" points="369" reactiontime="+96" swimtime="00:02:51.25" resultid="1924" heatid="6275" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:21.85" />
                    <SPLIT distance="150" swimtime="00:02:07.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="476" reactiontime="+96" swimtime="00:00:33.79" resultid="1925" heatid="6337" lane="2" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="2112">
              <RESULTS>
                <RESULT eventid="1198" points="535" reactiontime="+93" swimtime="00:02:54.78" resultid="2114" heatid="6115" lane="2" entrytime="00:02:53.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                    <SPLIT distance="100" swimtime="00:01:23.29" />
                    <SPLIT distance="150" swimtime="00:02:09.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="461" reactiontime="+88" swimtime="00:01:05.45" resultid="2115" heatid="6171" lane="1" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="543" reactiontime="+84" swimtime="00:00:34.66" resultid="2116" heatid="6214" lane="4" entrytime="00:00:34.37" />
                <RESULT eventid="1528" points="493" reactiontime="+83" swimtime="00:00:28.77" resultid="2117" heatid="6355" lane="2" entrytime="00:00:28.32" />
                <RESULT eventid="1610" points="541" reactiontime="+88" swimtime="00:01:17.53" resultid="2118" heatid="6405" lane="2" entrytime="00:01:18.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Delfin Inowrocław" nation="POL" region="KUJ">
          <CONTACT city="INOWROCŁAW" name="LEWANDOWSKI ZYGMUNT" street="WIERZBIŃSKIEGO" zip="88-100" />
          <ATHLETES>
            <ATHLETE birthdate="1937-09-19" firstname="ZYGMUNT" gender="M" lastname="LEWANDOWSKI" nation="POL" athleteid="1927">
              <RESULTS>
                <RESULT eventid="1137" points="634" swimtime="00:15:12.39" resultid="1928" heatid="6447" lane="4" entrytime="00:17:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.91" />
                    <SPLIT distance="100" swimtime="00:01:42.24" />
                    <SPLIT distance="200" swimtime="00:03:33.34" />
                    <SPLIT distance="300" swimtime="00:05:27.21" />
                    <SPLIT distance="400" swimtime="00:07:23.21" />
                    <SPLIT distance="500" swimtime="00:09:20.80" />
                    <SPLIT distance="600" swimtime="00:11:18.69" />
                    <SPLIT distance="700" swimtime="00:13:17.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="480" reactiontime="+89" swimtime="00:01:48.68" resultid="1929" heatid="6084" lane="1" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="367" reactiontime="+105" swimtime="00:00:50.27" resultid="1930" heatid="6225" lane="6" entrytime="00:00:50.00" entrycourse="SCM" />
                <RESULT eventid="1437" points="561" reactiontime="+99" swimtime="00:03:25.69" resultid="1931" heatid="6279" lane="1" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.85" />
                    <SPLIT distance="100" swimtime="00:01:36.36" />
                    <SPLIT distance="150" swimtime="00:02:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="444" reactiontime="+112" swimtime="00:02:00.65" resultid="1932" heatid="6317" lane="6" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="573" reactiontime="+111" swimtime="00:07:16.50" resultid="1933" heatid="6560" lane="3" entrytime="00:07:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.93" />
                    <SPLIT distance="100" swimtime="00:01:43.73" />
                    <SPLIT distance="150" swimtime="00:02:39.57" />
                    <SPLIT distance="200" swimtime="00:03:36.19" />
                    <SPLIT distance="250" swimtime="00:04:32.74" />
                    <SPLIT distance="300" swimtime="00:05:29.04" />
                    <SPLIT distance="350" swimtime="00:06:24.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Niezrzeszony Białystok" nation="POL">
          <CONTACT email="wzmasters@wp.pl" name="Żmiejko Wojciech" phone="797309140" />
          <ATHLETES>
            <ATHLETE birthdate="1963-01-01" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="1935">
              <RESULTS>
                <RESULT eventid="1168" points="783" reactiontime="+83" swimtime="00:01:08.99" resultid="1936" heatid="6096" lane="5" entrytime="00:01:09.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="746" reactiontime="+80" swimtime="00:01:00.37" resultid="1937" heatid="6174" lane="6" entrytime="00:01:00.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="761" reactiontime="+84" swimtime="00:00:29.99" resultid="1938" heatid="6235" lane="1" entrytime="00:00:30.25" />
                <RESULT eventid="1467" points="750" reactiontime="+85" swimtime="00:02:33.90" resultid="1939" heatid="6309" lane="1" entrytime="00:02:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:13.22" />
                    <SPLIT distance="150" swimtime="00:01:58.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="733" reactiontime="+87" swimtime="00:01:08.01" resultid="1940" heatid="6324" lane="1" entrytime="00:01:08.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="702" reactiontime="+82" swimtime="00:00:27.60" resultid="1941" heatid="6357" lane="3" entrytime="00:00:27.95" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Dęby Osielsko" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Adrian" gender="M" lastname="Teodorski" nation="POL" athleteid="2015">
              <RESULTS>
                <RESULT eventid="1092" points="538" reactiontime="+95" swimtime="00:05:24.62" resultid="2016" heatid="6492" lane="2" entrytime="00:05:18.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:06.65" />
                    <SPLIT distance="150" swimtime="00:01:48.97" />
                    <SPLIT distance="200" swimtime="00:02:31.02" />
                    <SPLIT distance="250" swimtime="00:03:19.75" />
                    <SPLIT distance="300" swimtime="00:04:10.79" />
                    <SPLIT distance="350" swimtime="00:04:48.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="705" reactiontime="+92" swimtime="00:01:06.50" resultid="2017" heatid="6100" lane="2" entrytime="00:01:02.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="621" reactiontime="+93" swimtime="00:00:57.85" resultid="2018" heatid="6179" lane="4" entrytime="00:00:56.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="718" reactiontime="+86" swimtime="00:00:27.70" resultid="2019" heatid="6239" lane="3" entrytime="00:00:27.80" />
                <RESULT eventid="1467" points="597" reactiontime="+92" swimtime="00:02:26.62" resultid="2020" heatid="6311" lane="6" entrytime="00:02:20.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:07.50" />
                    <SPLIT distance="150" swimtime="00:01:53.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="653" reactiontime="+91" swimtime="00:01:01.83" resultid="2021" heatid="6327" lane="5" entrytime="00:00:59.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="621" reactiontime="+77" swimtime="00:00:26.15" resultid="2022" heatid="6362" lane="6" entrytime="00:00:26.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="AZS UJ Kraków" nation="POL" region="KR">
          <CONTACT city="Kraków" name="Syryca Michał" phone="783-785-287" state="MAŁ" street="Piastowska 26 D" zip="30-065" />
          <ATHLETES>
            <ATHLETE birthdate="1992-08-01" firstname="Karolina" gender="F" lastname="Zadrożna" nation="POL" athleteid="2024">
              <RESULTS>
                <RESULT eventid="1122" points="535" swimtime="00:10:46.39" resultid="2025" heatid="6445" lane="3" entrytime="00:10:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:02:29.80" />
                    <SPLIT distance="200" swimtime="00:02:29.80" />
                    <SPLIT distance="400" swimtime="00:05:12.83" />
                    <SPLIT distance="500" swimtime="00:06:35.08" />
                    <SPLIT distance="600" swimtime="00:07:58.74" />
                    <SPLIT distance="700" swimtime="00:09:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="507" reactiontime="+59" swimtime="00:00:37.36" resultid="2026" heatid="6125" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1257" points="569" reactiontime="+92" swimtime="00:01:07.35" resultid="2027" heatid="6157" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="491" reactiontime="+61" swimtime="00:01:21.18" resultid="2028" heatid="6248" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="628" reactiontime="+92" swimtime="00:02:24.81" resultid="2029" heatid="6277" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:10.32" />
                    <SPLIT distance="150" swimtime="00:01:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="563" reactiontime="+87" swimtime="00:00:31.00" resultid="2030" heatid="6338" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1625" points="564" reactiontime="+91" swimtime="00:05:06.94" resultid="2031" heatid="6558" lane="2" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:12.98" />
                    <SPLIT distance="150" swimtime="00:01:52.05" />
                    <SPLIT distance="200" swimtime="00:02:31.38" />
                    <SPLIT distance="250" swimtime="00:03:10.83" />
                    <SPLIT distance="300" swimtime="00:03:50.44" />
                    <SPLIT distance="350" swimtime="00:04:30.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="BARAKUDA Legnica" nation="POL" region="DOL">
          <CONTACT email="jmalchar@o2.pl" name="Malchar Jowita" phone="506034671" />
          <ATHLETES>
            <ATHLETE birthdate="1982-12-28" firstname="Jowita" gender="F" lastname="Malchar" nation="POL" athleteid="2033">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. B" eventid="1058" points="508" reactiontime="+84" swimtime="00:06:14.78" resultid="2034" heatid="6431" lane="5" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:08.82" />
                    <SPLIT distance="200" swimtime="00:02:55.84" />
                    <SPLIT distance="250" swimtime="00:03:51.70" />
                    <SPLIT distance="300" swimtime="00:04:46.99" />
                    <SPLIT distance="350" swimtime="00:05:31.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="540" reactiontime="+82" swimtime="00:01:19.84" resultid="2035" heatid="6080" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="566" reactiontime="+81" swimtime="00:01:10.16" resultid="2036" heatid="6156" lane="6" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="503" reactiontime="+78" swimtime="00:00:41.82" resultid="2037" heatid="6198" lane="4" entrytime="00:00:44.00" />
                <RESULT eventid="1452" points="549" reactiontime="+78" swimtime="00:02:54.48" resultid="2038" heatid="6296" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                    <SPLIT distance="100" swimtime="00:01:22.35" />
                    <SPLIT distance="150" swimtime="00:02:13.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="502" reactiontime="+78" swimtime="00:01:29.80" resultid="2039" heatid="6508" lane="4" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="476" reactiontime="+76" swimtime="00:05:43.30" resultid="2040" heatid="6557" lane="5" entrytime="00:05:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:19.64" />
                    <SPLIT distance="150" swimtime="00:02:03.41" />
                    <SPLIT distance="200" swimtime="00:02:47.45" />
                    <SPLIT distance="250" swimtime="00:03:32.42" />
                    <SPLIT distance="300" swimtime="00:04:17.12" />
                    <SPLIT distance="350" swimtime="00:05:01.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-04-11" firstname="Sebastian" gender="M" lastname="Hudyka" nation="POL" athleteid="2041">
              <RESULTS>
                <RESULT eventid="1137" points="368" swimtime="00:12:01.88" resultid="2042" heatid="6451" lane="3" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                    <SPLIT distance="100" swimtime="00:01:27.37" />
                    <SPLIT distance="200" swimtime="00:03:00.08" />
                    <SPLIT distance="300" swimtime="00:04:31.72" />
                    <SPLIT distance="400" swimtime="00:06:04.97" />
                    <SPLIT distance="500" swimtime="00:07:38.74" />
                    <SPLIT distance="600" swimtime="00:09:12.84" />
                    <SPLIT distance="700" swimtime="00:10:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="374" reactiontime="+84" swimtime="00:01:14.08" resultid="2043" heatid="6165" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="386" reactiontime="+103" swimtime="00:02:42.57" resultid="2044" heatid="6283" lane="1" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:18.52" />
                    <SPLIT distance="150" swimtime="00:02:01.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="382" reactiontime="+95" swimtime="00:00:33.65" resultid="2045" heatid="6349" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1640" points="383" reactiontime="+97" swimtime="00:05:45.80" resultid="2046" heatid="6564" lane="4" entrytime="00:05:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                    <SPLIT distance="100" swimtime="00:01:23.14" />
                    <SPLIT distance="150" swimtime="00:02:07.99" />
                    <SPLIT distance="200" swimtime="00:02:52.56" />
                    <SPLIT distance="250" swimtime="00:03:36.81" />
                    <SPLIT distance="300" swimtime="00:04:21.01" />
                    <SPLIT distance="350" swimtime="00:05:04.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Start Poznań" nation="POL">
          <CONTACT city="Poznań" email="robert.beym@gmail.com" name="Beym Robert" phone="+48 512 111 513" street="Os. Batorego 8/67" zip="60-687" />
          <ATHLETES>
            <ATHLETE birthdate="1969-02-26" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="2048">
              <RESULTS>
                <RESULT eventid="1168" points="682" reactiontime="+80" swimtime="00:01:10.13" resultid="2049" heatid="6094" lane="1" entrytime="00:01:12.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="609" reactiontime="+77" swimtime="00:00:33.04" resultid="2050" heatid="6135" lane="1" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1393" points="617" reactiontime="+77" swimtime="00:01:11.33" resultid="2051" heatid="6259" lane="5" entrytime="00:01:11.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="629" reactiontime="+87" swimtime="00:02:39.11" resultid="2052" heatid="6307" lane="2" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:13.47" />
                    <SPLIT distance="150" swimtime="00:02:02.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="690" reactiontime="+76" swimtime="00:02:33.29" resultid="2053" heatid="6381" lane="6" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:52.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="508" reactiontime="+96" swimtime="00:05:14.83" resultid="2054" heatid="6565" lane="4" entrytime="00:05:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:01:55.00" />
                    <SPLIT distance="200" swimtime="00:02:35.72" />
                    <SPLIT distance="250" swimtime="00:03:15.93" />
                    <SPLIT distance="300" swimtime="00:03:55.89" />
                    <SPLIT distance="350" swimtime="00:04:35.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Rzeszów nizrzeszony" nation="POL" region="PDK" name.en="Rzeszow niezrzeszony">
          <CONTACT city="Rzeszów" email="wieslawcieklinski@wp.pl" name="Ciekliński" phone="602682904" state="PODKA" street="Jagiellońska 7/3" zip="35-025" />
          <ATHLETES>
            <ATHLETE birthdate="1957-06-08" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="2056">
              <RESULTS>
                <RESULT eventid="1168" points="470" reactiontime="+100" swimtime="00:01:27.46" resultid="2057" heatid="6087" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="602" reactiontime="+96" swimtime="00:01:09.49" resultid="2058" heatid="6166" lane="1" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="438" reactiontime="+74" swimtime="00:00:36.96" resultid="2059" heatid="6227" lane="5" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1437" points="554" reactiontime="+96" swimtime="00:02:40.43" resultid="2060" heatid="6282" lane="3" entrytime="00:02:44.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                    <SPLIT distance="150" swimtime="00:02:00.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="614" reactiontime="+86" swimtime="00:00:30.71" resultid="2061" heatid="6350" lane="4" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1640" points="538" reactiontime="+97" swimtime="00:05:51.88" resultid="2062" heatid="6563" lane="1" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:23.82" />
                    <SPLIT distance="150" swimtime="00:02:09.43" />
                    <SPLIT distance="200" swimtime="00:02:56.31" />
                    <SPLIT distance="250" swimtime="00:03:42.75" />
                    <SPLIT distance="300" swimtime="00:04:28.25" />
                    <SPLIT distance="350" swimtime="00:05:13.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="CityZen Masters Poznań" nation="POL" region="WIE">
          <CONTACT email="uks@ukscityzen.pl" internet="www.ukscityzen.pl" name="Roszak" />
          <ATHLETES>
            <ATHLETE birthdate="1988-01-01" firstname="Adrian" gender="M" lastname="Roszak" nation="POL" athleteid="2072">
              <RESULTS>
                <RESULT eventid="1137" points="616" swimtime="00:09:42.83" resultid="2073" heatid="6456" lane="6" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:08.21" />
                    <SPLIT distance="200" swimtime="00:02:19.54" />
                    <SPLIT distance="300" swimtime="00:03:31.96" />
                    <SPLIT distance="400" swimtime="00:04:45.19" />
                    <SPLIT distance="500" swimtime="00:05:59.28" />
                    <SPLIT distance="600" swimtime="00:07:14.46" />
                    <SPLIT distance="700" swimtime="00:08:30.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="750" reactiontime="+73" swimtime="00:00:54.34" resultid="2074" heatid="6180" lane="1" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="490" reactiontime="+93" swimtime="00:02:32.14" resultid="2075" heatid="6189" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:14.26" />
                    <SPLIT distance="150" swimtime="00:01:54.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="703" reactiontime="+72" swimtime="00:00:27.89" resultid="2076" heatid="6239" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1437" points="625" reactiontime="+76" swimtime="00:02:05.91" resultid="2077" heatid="6291" lane="2" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                    <SPLIT distance="100" swimtime="00:01:02.89" />
                    <SPLIT distance="150" swimtime="00:01:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="651" reactiontime="+77" swimtime="00:01:01.89" resultid="2078" heatid="6325" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="586" reactiontime="+94" swimtime="00:04:38.42" resultid="2079" heatid="6559" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:42.35" />
                    <SPLIT distance="200" swimtime="00:02:17.92" />
                    <SPLIT distance="250" swimtime="00:02:53.64" />
                    <SPLIT distance="300" swimtime="00:03:29.38" />
                    <SPLIT distance="350" swimtime="00:04:04.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Tadeusz" gender="M" lastname="Gołembiewski" nation="POL" athleteid="2080">
              <RESULTS>
                <RESULT eventid="1137" points="638" swimtime="00:09:45.52" resultid="2081" heatid="6456" lane="2" entrytime="00:09:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                    <SPLIT distance="200" swimtime="00:02:16.22" />
                    <SPLIT distance="300" swimtime="00:03:27.60" />
                    <SPLIT distance="400" swimtime="00:04:41.60" />
                    <SPLIT distance="500" swimtime="00:05:56.72" />
                    <SPLIT distance="600" swimtime="00:07:12.88" />
                    <SPLIT distance="700" swimtime="00:08:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="703" reactiontime="+81" swimtime="00:00:56.87" resultid="2082" heatid="6180" lane="6" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="622" reactiontime="+88" swimtime="00:02:27.45" resultid="2083" heatid="6190" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:10.03" />
                    <SPLIT distance="150" swimtime="00:01:48.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="691" reactiontime="+88" swimtime="00:00:28.68" resultid="2084" heatid="6240" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1437" points="674" reactiontime="+87" swimtime="00:02:06.20" resultid="2085" heatid="6291" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                    <SPLIT distance="100" swimtime="00:01:02.81" />
                    <SPLIT distance="150" swimtime="00:01:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="620" reactiontime="+83" swimtime="00:01:05.12" resultid="2086" heatid="6325" lane="3" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="682" reactiontime="+90" swimtime="00:04:34.26" resultid="2087" heatid="6560" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                    <SPLIT distance="100" swimtime="00:01:04.79" />
                    <SPLIT distance="150" swimtime="00:01:39.52" />
                    <SPLIT distance="200" swimtime="00:02:14.59" />
                    <SPLIT distance="250" swimtime="00:02:49.62" />
                    <SPLIT distance="300" swimtime="00:03:24.78" />
                    <SPLIT distance="350" swimtime="00:04:00.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Oświęcim" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1961-01-01" firstname="Tomasz" gender="M" lastname="Dorywalski" nation="POL" athleteid="2092">
              <RESULTS>
                <RESULT eventid="1228" points="609" reactiontime="+66" swimtime="00:00:36.11" resultid="2093" heatid="6133" lane="6" entrytime="00:00:36.50" />
                <RESULT eventid="1393" points="618" reactiontime="+65" swimtime="00:01:18.86" resultid="2094" heatid="6257" lane="6" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="630" reactiontime="+72" swimtime="00:02:53.68" resultid="2095" heatid="6377" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="100" swimtime="00:01:21.90" />
                    <SPLIT distance="150" swimtime="00:02:07.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="AZS UJCM Kraków" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1992-01-01" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" athleteid="2097">
              <RESULTS>
                <RESULT eventid="1153" points="905" reactiontime="+85" swimtime="00:01:09.26" resultid="2098" heatid="6082" lane="4" entrytime="00:01:08.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="703" reactiontime="+86" swimtime="00:02:50.88" resultid="2099" heatid="6107" lane="4" entrytime="00:02:46.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:21.85" />
                    <SPLIT distance="150" swimtime="00:02:06.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="751" swimtime="00:00:36.08" resultid="2100" heatid="6201" lane="2" entrytime="00:00:35.52" />
                <RESULT eventid="1452" points="768" reactiontime="+86" swimtime="00:02:31.70" resultid="2101" heatid="6298" lane="3" entrytime="00:02:26.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="743" reactiontime="+83" swimtime="00:00:28.27" resultid="2102" heatid="6340" lane="3" entrytime="00:00:27.62" />
                <RESULT eventid="1595" points="686" reactiontime="+87" swimtime="00:01:19.98" resultid="2103" heatid="6510" lane="4" entrytime="00:01:18.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UKS" name="UKS Trójka Oborniki" nation="POL" region="WIE">
          <CONTACT city="Oborniki" email="janwol@poczta.onet.pl" name="Wolniewicz Janusz" phone="791064667" state="WIE" street="Piłsudskiego 49/42" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-20" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" license="JanWol" athleteid="2120">
              <RESULTS>
                <RESULT eventid="1137" points="325" swimtime="00:14:42.96" resultid="2121" heatid="6448" lane="5" entrytime="00:14:43.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:38.84" />
                    <SPLIT distance="200" swimtime="00:03:25.43" />
                    <SPLIT distance="300" swimtime="00:05:14.03" />
                    <SPLIT distance="400" swimtime="00:07:05.66" />
                    <SPLIT distance="500" swimtime="00:08:59.24" />
                    <SPLIT distance="600" swimtime="00:10:55.00" />
                    <SPLIT distance="700" swimtime="00:12:51.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="450" reactiontime="+101" swimtime="00:01:21.34" resultid="2122" heatid="6162" lane="5" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="389" swimtime="00:03:13.30" resultid="2123" heatid="6280" lane="2" entrytime="00:03:09.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:01:33.31" />
                    <SPLIT distance="150" swimtime="00:02:24.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="444" reactiontime="+101" swimtime="00:00:35.77" resultid="2124" heatid="6345" lane="5" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1640" points="329" reactiontime="+107" swimtime="00:07:07.05" resultid="2125" heatid="6561" lane="4" entrytime="00:06:50.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.01" />
                    <SPLIT distance="100" swimtime="00:01:41.65" />
                    <SPLIT distance="150" swimtime="00:02:36.04" />
                    <SPLIT distance="200" swimtime="00:03:31.24" />
                    <SPLIT distance="250" swimtime="00:04:25.74" />
                    <SPLIT distance="300" swimtime="00:05:20.15" />
                    <SPLIT distance="350" swimtime="00:06:12.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KOROKRAK" name="Masters Korona Kraków" nation="POL" region="KR">
          <CONTACT email="masterskorona@wp.pl" internet="www.masterskorona.pl" name="Mariola Kuliś" phone="500677133" state="MAŁ" street="Kalwaryjska" />
          <ATHLETES>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="2129">
              <RESULTS>
                <RESULT eventid="1153" points="776" reactiontime="+74" swimtime="00:01:18.04" resultid="2130" heatid="6077" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="781" reactiontime="+67" swimtime="00:00:36.23" resultid="2131" heatid="6120" lane="3" entrytime="00:00:50.50" />
                <RESULT eventid="1318" points="761" reactiontime="+78" swimtime="00:00:39.51" resultid="2132" heatid="6196" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1378" points="738" reactiontime="+68" swimtime="00:01:20.89" resultid="2133" heatid="6248" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="704" reactiontime="+72" swimtime="00:00:31.65" resultid="2134" heatid="6332" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1543" points="742" reactiontime="+67" swimtime="00:02:59.32" resultid="2135" heatid="6368" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                    <SPLIT distance="100" swimtime="00:01:27.40" />
                    <SPLIT distance="150" swimtime="00:02:14.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="2136">
              <RESULTS>
                <RESULT eventid="1257" points="620" reactiontime="+95" swimtime="00:01:14.49" resultid="2137" heatid="6156" lane="1" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="650" reactiontime="+79" swimtime="00:00:35.20" resultid="2138" heatid="6222" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1452" points="706" reactiontime="+85" swimtime="00:02:58.61" resultid="2139" heatid="6297" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:23.93" />
                    <SPLIT distance="150" swimtime="00:02:16.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="660" reactiontime="+89" swimtime="00:01:20.82" resultid="2140" heatid="6315" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-26" firstname="Marta" gender="F" lastname="Wysocka" nation="POL" athleteid="2141">
              <RESULTS>
                <RESULT eventid="1183" points="730" reactiontime="+93" swimtime="00:03:18.21" resultid="2142" heatid="6106" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.71" />
                    <SPLIT distance="100" swimtime="00:01:32.75" />
                    <SPLIT distance="150" swimtime="00:02:25.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="739" reactiontime="+84" swimtime="00:00:41.92" resultid="2143" heatid="6199" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1595" points="788" reactiontime="+85" swimtime="00:01:30.23" resultid="2144" heatid="6509" lane="2" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-22" firstname="Alicja" gender="F" lastname="Romańska" nation="POL" athleteid="2145">
              <RESULTS>
                <RESULT eventid="1122" points="228" swimtime="00:15:15.89" resultid="2146" heatid="6442" lane="5" entrytime="00:15:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.88" />
                    <SPLIT distance="200" swimtime="00:03:47.78" />
                    <SPLIT distance="300" swimtime="00:05:43.15" />
                    <SPLIT distance="400" swimtime="00:07:39.36" />
                    <SPLIT distance="500" swimtime="00:09:34.40" />
                    <SPLIT distance="600" swimtime="00:11:27.14" />
                    <SPLIT distance="700" swimtime="00:13:21.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" status="DNS" swimtime="00:00:00.00" resultid="2147" heatid="6076" lane="6" entrytime="00:01:50.00" />
                <RESULT eventid="1257" points="199" reactiontime="+101" swimtime="00:01:38.73" resultid="2148" heatid="6150" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="129" reactiontime="+113" swimtime="00:00:57.80" resultid="2149" heatid="6218" lane="3" entrytime="00:00:58.01" />
                <RESULT eventid="1422" points="204" reactiontime="+114" swimtime="00:03:33.45" resultid="2150" heatid="6272" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.34" />
                    <SPLIT distance="100" swimtime="00:01:44.31" />
                    <SPLIT distance="150" swimtime="00:02:40.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" reactiontime="+109" status="DNS" swimtime="00:00:00.00" resultid="2151" heatid="6312" lane="2" entrytime="00:02:05.00" />
                <RESULT eventid="1513" points="228" reactiontime="+99" swimtime="00:00:43.81" resultid="2152" heatid="6331" lane="2" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-07-26" firstname="Anna" gender="F" lastname="Kożmin" nation="POL" athleteid="2153">
              <RESULTS>
                <RESULT eventid="1153" points="360" reactiontime="+119" swimtime="00:01:55.27" resultid="2154" heatid="6074" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="331" reactiontime="+115" swimtime="00:04:30.15" resultid="2155" heatid="6103" lane="2" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.82" />
                    <SPLIT distance="100" swimtime="00:02:06.81" />
                    <SPLIT distance="150" swimtime="00:03:19.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="415" swimtime="00:00:51.73" resultid="2156" heatid="6195" lane="2" entrytime="00:00:53.00" />
                <RESULT eventid="1452" points="320" reactiontime="+112" swimtime="00:04:23.30" resultid="2157" heatid="6293" lane="4" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.57" />
                    <SPLIT distance="100" swimtime="00:02:07.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="371" reactiontime="+108" swimtime="00:02:00.28" resultid="2158" heatid="6505" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-15" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="2159">
              <RESULTS>
                <RESULT eventid="1153" points="233" reactiontime="+105" swimtime="00:02:27.77" resultid="2160" heatid="6074" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="284" reactiontime="+119" swimtime="00:05:28.85" resultid="2161" heatid="6102" lane="4" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.55" />
                    <SPLIT distance="100" swimtime="00:02:36.96" />
                    <SPLIT distance="150" swimtime="00:04:05.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="131" reactiontime="+118" swimtime="00:01:17.21" resultid="2162" heatid="6218" lane="5" entrytime="00:01:22.00" />
                <RESULT eventid="1422" points="189" reactiontime="+126" swimtime="00:04:55.33" resultid="2163" heatid="6271" lane="6" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.86" />
                    <SPLIT distance="100" swimtime="00:02:10.67" />
                    <SPLIT distance="150" swimtime="00:03:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="212" reactiontime="+110" swimtime="00:00:58.32" resultid="2164" heatid="6330" lane="1" entrytime="00:00:59.00" />
                <RESULT eventid="1595" points="316" reactiontime="+118" swimtime="00:02:22.64" resultid="2165" heatid="6504" lane="4" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-04-24" firstname="Krzysztof" gender="M" lastname="Chołda" nation="POL" athleteid="2166">
              <RESULTS>
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="2167" heatid="6451" lane="5" entrytime="00:12:08.00" />
                <RESULT eventid="1168" points="427" reactiontime="+94" swimtime="00:01:24.43" resultid="2168" heatid="6089" lane="1" entrytime="00:01:24.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="2169" heatid="6166" lane="5" entrytime="00:01:10.56" />
                <RESULT eventid="1333" points="418" reactiontime="+91" swimtime="00:00:41.07" resultid="2170" heatid="6209" lane="5" entrytime="00:00:41.55" />
                <RESULT eventid="1467" points="406" reactiontime="+93" swimtime="00:03:08.70" resultid="2171" heatid="6304" lane="6" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:31.79" />
                    <SPLIT distance="150" swimtime="00:02:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="479" reactiontime="+89" swimtime="00:00:31.35" resultid="2172" heatid="6350" lane="5" entrytime="00:00:31.14" />
                <RESULT eventid="1610" points="402" reactiontime="+91" swimtime="00:01:33.15" resultid="2173" heatid="6400" lane="6" entrytime="00:01:34.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-04" firstname="Andrzej" gender="M" lastname="Data" nation="POL" athleteid="2174">
              <RESULTS>
                <RESULT eventid="1137" points="367" swimtime="00:13:11.64" resultid="2175" heatid="6450" lane="4" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:23.64" />
                    <SPLIT distance="200" swimtime="00:03:01.11" />
                    <SPLIT distance="300" swimtime="00:04:42.08" />
                    <SPLIT distance="400" swimtime="00:06:24.70" />
                    <SPLIT distance="500" swimtime="00:08:13.47" />
                    <SPLIT distance="600" swimtime="00:09:52.45" />
                    <SPLIT distance="700" swimtime="00:11:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="419" reactiontime="+99" swimtime="00:03:35.40" resultid="2176" heatid="6112" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                    <SPLIT distance="100" swimtime="00:01:41.10" />
                    <SPLIT distance="150" swimtime="00:02:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="404" reactiontime="+96" swimtime="00:01:16.93" resultid="2177" heatid="6163" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="351" reactiontime="+124" swimtime="00:00:45.63" resultid="2178" heatid="6207" lane="1" entrytime="00:00:44.00" />
                <RESULT eventid="1437" points="352" reactiontime="+94" swimtime="00:02:56.01" resultid="2179" heatid="6284" lane="6" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:20.94" />
                    <SPLIT distance="150" swimtime="00:02:08.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="411" reactiontime="+97" swimtime="00:01:37.82" resultid="2180" heatid="6399" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="363" reactiontime="+109" swimtime="00:06:16.17" resultid="2181" heatid="6563" lane="6" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                    <SPLIT distance="100" swimtime="00:01:21.06" />
                    <SPLIT distance="150" swimtime="00:02:07.86" />
                    <SPLIT distance="200" swimtime="00:02:56.45" />
                    <SPLIT distance="250" swimtime="00:03:47.35" />
                    <SPLIT distance="300" swimtime="00:04:38.08" />
                    <SPLIT distance="350" swimtime="00:05:28.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-03-07" firstname="Robert" gender="M" lastname="Grela" nation="POL" athleteid="2182">
              <RESULTS>
                <RESULT eventid="1363" points="698" reactiontime="+79" swimtime="00:00:30.05" resultid="2183" heatid="6238" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1498" points="641" reactiontime="+79" swimtime="00:01:08.03" resultid="2184" heatid="6325" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-15" firstname="Michał" gender="M" lastname="Gugała" nation="POL" athleteid="2185">
              <RESULTS>
                <RESULT eventid="1137" points="289" swimtime="00:12:33.46" resultid="2186" heatid="6449" lane="4" entrytime="00:13:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="200" swimtime="00:02:54.38" />
                    <SPLIT distance="300" swimtime="00:04:29.91" />
                    <SPLIT distance="400" swimtime="00:07:05.40" />
                    <SPLIT distance="500" swimtime="00:07:42.14" />
                    <SPLIT distance="600" swimtime="00:09:20.53" />
                    <SPLIT distance="700" swimtime="00:10:59.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="411" reactiontime="+108" swimtime="00:01:08.12" resultid="2187" heatid="6163" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="306" reactiontime="+105" swimtime="00:05:56.88" resultid="2188" heatid="6562" lane="4" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:13.34" />
                    <SPLIT distance="150" swimtime="00:01:57.49" />
                    <SPLIT distance="200" swimtime="00:02:45.15" />
                    <SPLIT distance="250" swimtime="00:03:32.99" />
                    <SPLIT distance="300" swimtime="00:04:22.29" />
                    <SPLIT distance="350" swimtime="00:05:11.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-15" firstname="Mariusz" gender="M" lastname="Kaliszyk" nation="POL" athleteid="2189">
              <RESULTS>
                <RESULT eventid="1272" points="709" reactiontime="+78" swimtime="00:00:59.89" resultid="2190" heatid="6167" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="739" reactiontime="+77" swimtime="00:00:29.48" resultid="2191" heatid="6229" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1528" points="707" reactiontime="+78" swimtime="00:00:27.40" resultid="2192" heatid="6349" lane="2" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-26" firstname="Anna" gender="F" lastname="Kasprzykowska" nation="POL" athleteid="2193">
              <RESULTS>
                <RESULT eventid="1348" points="159" swimtime="00:00:53.20" resultid="2194" heatid="6218" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1422" points="156" reactiontime="+97" swimtime="00:03:52.72" resultid="2195" heatid="6271" lane="3" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.40" />
                    <SPLIT distance="100" swimtime="00:01:51.34" />
                    <SPLIT distance="150" swimtime="00:02:52.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-05-16" firstname="Tadeusz" gender="M" lastname="Krawczyk" nation="POL" athleteid="2196">
              <RESULTS>
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="2197" heatid="6446" lane="2" />
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="2198" heatid="6083" lane="2" entrytime="00:02:15.00" />
                <RESULT eventid="1228" points="154" reactiontime="+72" swimtime="00:01:05.76" resultid="2199" heatid="6127" lane="1" entrytime="00:00:58.00" />
                <RESULT eventid="1393" reactiontime="+99" status="DSQ" swimtime="00:02:26.74" resultid="2200" heatid="6251" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="2201" heatid="6280" lane="6" entrytime="00:03:20.00" />
                <RESULT eventid="1528" points="254" reactiontime="+111" swimtime="00:00:44.60" resultid="2202" heatid="6343" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-06-03" firstname="Antoni" gender="M" lastname="Kubis" nation="POL" athleteid="2203">
              <RESULTS>
                <RESULT eventid="1168" points="388" reactiontime="+123" swimtime="00:01:43.56" resultid="2204" heatid="6085" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="318" reactiontime="+113" swimtime="00:00:46.64" resultid="2205" heatid="6224" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1528" points="243" reactiontime="+132" swimtime="00:00:45.26" resultid="2206" heatid="6342" lane="3" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-10-12" firstname="Joanna" gender="F" lastname="Kwatera" nation="POL" athleteid="2207">
              <RESULTS>
                <RESULT eventid="1183" points="509" reactiontime="+82" swimtime="00:03:17.61" resultid="2208" heatid="6106" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.57" />
                    <SPLIT distance="100" swimtime="00:01:32.66" />
                    <SPLIT distance="150" swimtime="00:02:24.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="521" reactiontime="+82" swimtime="00:00:42.35" resultid="2209" heatid="6199" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1595" points="436" reactiontime="+77" swimtime="00:01:33.19" resultid="2210" heatid="6509" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-16" firstname="Kamil" gender="M" lastname="Latuszek" nation="POL" athleteid="2211">
              <RESULTS>
                <RESULT eventid="1168" points="622" reactiontime="+77" swimtime="00:01:09.32" resultid="2212" heatid="6095" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="579" reactiontime="+75" swimtime="00:00:59.22" resultid="2213" heatid="6177" lane="3" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="493" reactiontime="+76" swimtime="00:02:16.25" resultid="2214" heatid="6288" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:06.58" />
                    <SPLIT distance="150" swimtime="00:01:42.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="602" reactiontime="+73" swimtime="00:00:26.43" resultid="2215" heatid="6361" lane="1" entrytime="00:00:26.70" />
                <RESULT eventid="1640" points="440" reactiontime="+76" swimtime="00:05:06.26" resultid="2216" heatid="6569" lane="3" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                    <SPLIT distance="150" swimtime="00:01:46.46" />
                    <SPLIT distance="200" swimtime="00:02:25.15" />
                    <SPLIT distance="250" swimtime="00:03:04.09" />
                    <SPLIT distance="300" swimtime="00:03:44.08" />
                    <SPLIT distance="350" swimtime="00:04:24.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="2217">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. G" eventid="1058" points="580" reactiontime="+109" swimtime="00:07:23.34" resultid="2218" heatid="6430" lane="1" entrytime="00:07:32.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.42" />
                    <SPLIT distance="100" swimtime="00:01:47.52" />
                    <SPLIT distance="150" swimtime="00:02:44.11" />
                    <SPLIT distance="200" swimtime="00:03:39.97" />
                    <SPLIT distance="250" swimtime="00:04:41.38" />
                    <SPLIT distance="300" swimtime="00:05:43.80" />
                    <SPLIT distance="350" swimtime="00:06:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="564" reactiontime="+104" swimtime="00:01:33.74" resultid="2219" heatid="6078" lane="1" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. G" eventid="1287" points="545" reactiontime="+122" swimtime="00:03:47.51" resultid="2220" heatid="6182" lane="5" entrytime="00:03:49.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.89" />
                    <SPLIT distance="100" swimtime="00:01:50.03" />
                    <SPLIT distance="150" swimtime="00:02:49.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="531" reactiontime="+102" swimtime="00:00:41.44" resultid="2221" heatid="6220" lane="6" entrytime="00:00:43.01" />
                <RESULT eventid="1452" points="548" reactiontime="+113" swimtime="00:03:30.77" resultid="2222" heatid="6295" lane="6" entrytime="00:03:34.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.03" />
                    <SPLIT distance="100" swimtime="00:01:44.21" />
                    <SPLIT distance="150" swimtime="00:02:44.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="410" reactiontime="+110" swimtime="00:01:43.76" resultid="2223" heatid="6313" lane="4" entrytime="00:01:41.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="565" reactiontime="+110" swimtime="00:06:43.39" resultid="2224" heatid="6554" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                    <SPLIT distance="100" swimtime="00:01:35.14" />
                    <SPLIT distance="150" swimtime="00:02:28.18" />
                    <SPLIT distance="200" swimtime="00:03:20.44" />
                    <SPLIT distance="250" swimtime="00:04:12.55" />
                    <SPLIT distance="300" swimtime="00:05:03.08" />
                    <SPLIT distance="350" swimtime="00:05:54.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-17" firstname="Wojciech" gender="M" lastname="Liszkowski" nation="POL" athleteid="2225">
              <RESULTS>
                <RESULT eventid="1333" points="598" swimtime="00:00:35.00" resultid="2226" heatid="6210" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1363" points="752" reactiontime="+81" swimtime="00:00:29.31" resultid="2227" heatid="6233" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1610" points="611" reactiontime="+76" swimtime="00:01:19.16" resultid="2228" heatid="6401" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="2229">
              <RESULTS>
                <RESULT eventid="1137" points="567" swimtime="00:13:40.76" resultid="2230" heatid="6448" lane="4" entrytime="00:14:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:36.45" />
                    <SPLIT distance="200" swimtime="00:03:20.76" />
                    <SPLIT distance="300" swimtime="00:05:05.48" />
                    <SPLIT distance="400" swimtime="00:06:49.04" />
                    <SPLIT distance="500" swimtime="00:08:33.13" />
                    <SPLIT distance="600" swimtime="00:10:15.80" />
                    <SPLIT distance="700" swimtime="00:11:58.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="771" reactiontime="+120" swimtime="00:01:11.99" resultid="2231" heatid="6165" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="415" reactiontime="+130" swimtime="00:04:05.98" resultid="2232" heatid="6185" lane="5" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.34" />
                    <SPLIT distance="100" swimtime="00:02:00.87" />
                    <SPLIT distance="150" swimtime="00:03:06.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="634" reactiontime="+119" swimtime="00:02:52.98" resultid="2233" heatid="6281" lane="2" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:01:20.44" />
                    <SPLIT distance="150" swimtime="00:02:07.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="474" reactiontime="+125" swimtime="00:03:41.72" resultid="2234" heatid="6302" lane="1" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.64" />
                    <SPLIT distance="100" swimtime="00:01:52.25" />
                    <SPLIT distance="150" swimtime="00:02:56.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="667" reactiontime="+106" swimtime="00:00:32.35" resultid="2235" heatid="6347" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1640" points="634" reactiontime="+135" swimtime="00:06:20.75" resultid="2236" heatid="6562" lane="1" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.90" />
                    <SPLIT distance="100" swimtime="00:01:33.46" />
                    <SPLIT distance="150" swimtime="00:02:21.62" />
                    <SPLIT distance="200" swimtime="00:03:11.04" />
                    <SPLIT distance="250" swimtime="00:04:00.71" />
                    <SPLIT distance="300" swimtime="00:04:49.43" />
                    <SPLIT distance="350" swimtime="00:05:37.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-01" firstname="Paulina" gender="F" lastname="Palmowska" nation="POL" athleteid="2237">
              <RESULTS>
                <RESULT eventid="1213" points="685" reactiontime="+65" swimtime="00:00:34.54" resultid="2238" heatid="6125" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1257" points="572" reactiontime="+71" swimtime="00:01:09.22" resultid="2239" heatid="6158" lane="2" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="604" reactiontime="+73" swimtime="00:01:15.07" resultid="2240" heatid="6248" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="519" reactiontime="+73" swimtime="00:02:56.57" resultid="2241" heatid="6298" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:21.20" />
                    <SPLIT distance="150" swimtime="00:02:12.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="522" reactiontime="+70" swimtime="00:02:47.83" resultid="2242" heatid="6371" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                    <SPLIT distance="100" swimtime="00:01:19.72" />
                    <SPLIT distance="150" swimtime="00:02:03.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="463" reactiontime="+77" swimtime="00:05:43.73" resultid="2243" heatid="6558" lane="6" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                    <SPLIT distance="100" swimtime="00:01:24.92" />
                    <SPLIT distance="150" swimtime="00:02:08.49" />
                    <SPLIT distance="200" swimtime="00:02:52.15" />
                    <SPLIT distance="250" swimtime="00:03:36.20" />
                    <SPLIT distance="300" swimtime="00:04:20.03" />
                    <SPLIT distance="350" swimtime="00:05:03.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="2244">
              <RESULTS>
                <RESULT eventid="1168" points="624" reactiontime="+90" swimtime="00:01:16.67" resultid="2245" heatid="6092" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="669" reactiontime="+77" swimtime="00:00:35.01" resultid="2246" heatid="6133" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1363" points="686" reactiontime="+94" swimtime="00:00:31.43" resultid="2247" heatid="6231" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1393" status="DNS" swimtime="00:00:00.00" resultid="2248" heatid="6257" lane="4" entrytime="00:01:16.00" />
                <RESULT eventid="1498" points="586" reactiontime="+91" swimtime="00:01:15.46" resultid="2249" heatid="6322" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="2250" heatid="6378" lane="4" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-18" firstname="Bartosz" gender="M" lastname="Próchniewicz" nation="POL" athleteid="2251">
              <RESULTS>
                <RESULT eventid="1228" points="124" reactiontime="+69" swimtime="00:00:52.26" resultid="2252" heatid="6128" lane="6" entrytime="00:00:52.83" />
                <RESULT eventid="1393" points="112" reactiontime="+73" swimtime="00:01:57.30" resultid="2253" heatid="6252" lane="4" entrytime="00:01:40.00" />
                <RESULT eventid="1528" points="110" reactiontime="+83" swimtime="00:00:48.02" resultid="2254" heatid="6343" lane="1" entrytime="00:00:43.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-12-18" firstname="Szymon" gender="M" lastname="Pyrć" nation="POL" athleteid="2255">
              <RESULTS>
                <RESULT eventid="1137" points="578" swimtime="00:10:18.37" resultid="2256" heatid="6452" lane="1" entrytime="00:11:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:13.18" />
                    <SPLIT distance="200" swimtime="00:02:30.71" />
                    <SPLIT distance="300" swimtime="00:03:48.69" />
                    <SPLIT distance="400" swimtime="00:05:07.00" />
                    <SPLIT distance="500" swimtime="00:06:25.24" />
                    <SPLIT distance="600" swimtime="00:07:43.27" />
                    <SPLIT distance="700" swimtime="00:09:01.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="628" reactiontime="+83" swimtime="00:02:31.61" resultid="2257" heatid="6190" lane="2" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:12.36" />
                    <SPLIT distance="150" swimtime="00:01:52.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="510" reactiontime="+84" swimtime="00:00:31.46" resultid="2258" heatid="6236" lane="1" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="2259">
              <RESULTS>
                <RESULT eventid="1183" points="204" reactiontime="+120" swimtime="00:04:37.35" resultid="2260" heatid="6102" lane="3" entrytime="00:04:36.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.96" />
                    <SPLIT distance="100" swimtime="00:02:14.83" />
                    <SPLIT distance="150" swimtime="00:03:25.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="166" reactiontime="+80" swimtime="00:00:57.14" resultid="2261" heatid="6120" lane="1" entrytime="00:00:55.32" />
                <RESULT eventid="1318" points="184" reactiontime="+118" swimtime="00:00:59.71" resultid="2262" heatid="6194" lane="1" entrytime="00:00:57.96" />
                <RESULT eventid="1378" points="137" reactiontime="+64" swimtime="00:02:09.11" resultid="2263" heatid="6244" lane="6" entrytime="00:02:05.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="2264" heatid="6367" lane="2" entrytime="00:04:33.63" />
                <RESULT eventid="1595" points="190" reactiontime="+117" swimtime="00:02:10.63" resultid="2265" heatid="6504" lane="2" entrytime="00:02:12.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-28" firstname="Wojciech" gender="M" lastname="Wolski" nation="POL" athleteid="2266">
              <RESULTS>
                <RESULT eventid="1528" points="439" reactiontime="+91" swimtime="00:00:32.26" resultid="2267" heatid="6348" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1610" points="499" reactiontime="+83" swimtime="00:01:26.66" resultid="2268" heatid="6402" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-12-07" firstname="Jarosław" gender="M" lastname="Zadrożny" nation="POL" athleteid="2269">
              <RESULTS>
                <RESULT eventid="1137" points="407" swimtime="00:12:22.14" resultid="2270" heatid="6450" lane="2" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                    <SPLIT distance="100" swimtime="00:01:24.68" />
                    <SPLIT distance="200" swimtime="00:02:56.28" />
                    <SPLIT distance="300" swimtime="00:04:28.55" />
                    <SPLIT distance="400" swimtime="00:06:02.28" />
                    <SPLIT distance="500" swimtime="00:07:39.34" />
                    <SPLIT distance="600" swimtime="00:09:15.12" />
                    <SPLIT distance="700" swimtime="00:10:51.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="446" swimtime="00:01:11.65" resultid="2271" heatid="6164" lane="2" entrytime="00:01:13.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" status="DNS" swimtime="00:00:00.00" resultid="2272" heatid="6228" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1437" points="422" reactiontime="+86" swimtime="00:02:43.32" resultid="2273" heatid="6281" lane="4" entrytime="00:02:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                    <SPLIT distance="150" swimtime="00:02:01.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="431" reactiontime="+85" swimtime="00:00:32.47" resultid="2274" heatid="6347" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1640" points="421" reactiontime="+93" swimtime="00:05:50.34" resultid="2275" heatid="6563" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:20.17" />
                    <SPLIT distance="150" swimtime="00:02:04.11" />
                    <SPLIT distance="200" swimtime="00:02:48.81" />
                    <SPLIT distance="250" swimtime="00:03:34.05" />
                    <SPLIT distance="300" swimtime="00:04:19.96" />
                    <SPLIT distance="350" swimtime="00:05:06.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-07" firstname="Sandra" gender="F" lastname="Pęczek" nation="POL" athleteid="2276">
              <RESULTS>
                <RESULT eventid="1153" points="622" reactiontime="+84" swimtime="00:01:16.83" resultid="2277" heatid="6082" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" status="DNS" swimtime="00:00:00.00" resultid="2278" heatid="6158" lane="5" entrytime="00:01:07.00" />
                <RESULT eventid="1318" points="814" reactiontime="+78" swimtime="00:00:36.51" resultid="2279" heatid="6201" lane="5" entrytime="00:00:36.50" />
                <RESULT eventid="1595" points="578" reactiontime="+82" swimtime="00:01:24.88" resultid="2280" heatid="6510" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-27" firstname="Wacław" gender="M" lastname="Brożek" nation="POL" athleteid="2281">
              <RESULTS>
                <RESULT eventid="1137" points="279" swimtime="00:14:01.58" resultid="2282" heatid="6449" lane="5" entrytime="00:13:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.34" />
                    <SPLIT distance="200" swimtime="00:03:17.49" />
                    <SPLIT distance="300" swimtime="00:05:03.98" />
                    <SPLIT distance="400" swimtime="00:06:50.98" />
                    <SPLIT distance="500" swimtime="00:08:39.64" />
                    <SPLIT distance="600" swimtime="00:10:29.04" />
                    <SPLIT distance="700" swimtime="00:12:14.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="303" reactiontime="+92" swimtime="00:01:34.64" resultid="2283" heatid="6085" lane="4" entrytime="00:01:38.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="182" reactiontime="+90" swimtime="00:00:50.90" resultid="2284" heatid="6127" lane="4" entrytime="00:00:56.00" />
                <RESULT eventid="1363" points="323" reactiontime="+111" swimtime="00:00:39.90" resultid="2285" heatid="6224" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1467" points="279" reactiontime="+98" swimtime="00:03:33.84" resultid="2286" heatid="6302" lane="5" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:01:42.00" />
                    <SPLIT distance="150" swimtime="00:02:46.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="295" reactiontime="+90" swimtime="00:06:34.35" resultid="2287" heatid="6562" lane="6" entrytime="00:06:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                    <SPLIT distance="100" swimtime="00:01:33.37" />
                    <SPLIT distance="150" swimtime="00:02:21.87" />
                    <SPLIT distance="200" swimtime="00:03:10.42" />
                    <SPLIT distance="250" swimtime="00:04:01.46" />
                    <SPLIT distance="300" swimtime="00:04:53.09" />
                    <SPLIT distance="350" swimtime="00:05:45.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-08-25" firstname="Mieczysław" gender="M" lastname="Strąk" nation="POL" athleteid="2288">
              <RESULTS>
                <RESULT eventid="1333" points="201" reactiontime="+114" swimtime="00:00:56.61" resultid="2289" heatid="6203" lane="6" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="2290">
              <RESULTS>
                <RESULT eventid="1058" points="390" reactiontime="+99" swimtime="00:07:15.56" resultid="2291" heatid="6430" lane="5" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.45" />
                    <SPLIT distance="100" swimtime="00:01:51.08" />
                    <SPLIT distance="150" swimtime="00:02:45.37" />
                    <SPLIT distance="200" swimtime="00:03:39.36" />
                    <SPLIT distance="250" swimtime="00:04:39.56" />
                    <SPLIT distance="300" swimtime="00:05:38.28" />
                    <SPLIT distance="350" swimtime="00:06:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="424" reactiontime="+91" swimtime="00:01:31.02" resultid="2292" heatid="6077" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="419" reactiontime="+80" swimtime="00:00:42.00" resultid="2293" heatid="6121" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1378" points="372" reactiontime="+87" swimtime="00:01:32.70" resultid="2294" heatid="6245" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="370" reactiontime="+93" swimtime="00:03:25.84" resultid="2295" heatid="6294" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.91" />
                    <SPLIT distance="100" swimtime="00:01:37.79" />
                    <SPLIT distance="150" swimtime="00:02:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="405" reactiontime="+88" swimtime="00:03:16.54" resultid="2296" heatid="6368" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:37.30" />
                    <SPLIT distance="150" swimtime="00:02:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="332" reactiontime="+106" swimtime="00:06:32.58" resultid="2297" heatid="6556" lane="5" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                    <SPLIT distance="100" swimtime="00:01:28.15" />
                    <SPLIT distance="150" swimtime="00:02:17.04" />
                    <SPLIT distance="200" swimtime="00:03:08.40" />
                    <SPLIT distance="250" swimtime="00:04:00.28" />
                    <SPLIT distance="300" swimtime="00:04:52.52" />
                    <SPLIT distance="350" swimtime="00:05:44.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-06-20" firstname="Tomasz" gender="M" lastname="Kalawa" nation="POL" athleteid="2298">
              <RESULTS>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="2299" heatid="6347" lane="5" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-03-21" firstname="Janusz" gender="M" lastname="Gołębiewski" nation="POL" athleteid="2300">
              <RESULTS>
                <RESULT eventid="1198" points="98" swimtime="00:06:22.13" resultid="2301" heatid="6109" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.00" />
                    <SPLIT distance="100" swimtime="00:02:57.81" />
                    <SPLIT distance="150" swimtime="00:04:41.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="172" reactiontime="+161" swimtime="00:01:01.50" resultid="2302" heatid="6202" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1610" points="129" reactiontime="+139" swimtime="00:02:36.04" resultid="2303" heatid="6396" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-15" firstname="Monika" gender="F" lastname="Jaworska" nation="POL" athleteid="2304">
              <RESULTS>
                <RESULT eventid="1348" points="545" reactiontime="+85" swimtime="00:00:33.77" resultid="2305" heatid="6222" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1513" points="516" reactiontime="+85" swimtime="00:00:31.92" resultid="2306" heatid="6339" lane="6" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-08" firstname="Tomasz" gender="M" lastname="Czerniecki" nation="POL" athleteid="2307">
              <RESULTS>
                <RESULT eventid="1528" points="650" reactiontime="+74" swimtime="00:00:26.63" resultid="2308" heatid="6363" lane="2" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-10-18" firstname="Dorota" gender="F" lastname="WIDZ-SZWARC" nation="POL" athleteid="2309">
              <RESULTS>
                <RESULT eventid="1257" points="420" reactiontime="+105" swimtime="00:01:24.81" resultid="2310" heatid="6154" lane="5" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="378" reactiontime="+106" swimtime="00:03:10.67" resultid="2311" heatid="6275" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                    <SPLIT distance="100" swimtime="00:01:28.48" />
                    <SPLIT distance="150" swimtime="00:02:19.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="429" reactiontime="+105" swimtime="00:00:37.32" resultid="2312" heatid="6334" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-24" firstname="Robert" gender="M" lastname="Trzos" nation="POL" athleteid="2314">
              <RESULTS>
                <RESULT eventid="1198" points="527" reactiontime="+82" swimtime="00:02:55.50" resultid="2315" heatid="6114" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                    <SPLIT distance="150" swimtime="00:02:09.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="430" reactiontime="+81" swimtime="00:00:38.17" resultid="2316" heatid="6211" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1610" points="433" reactiontime="+78" swimtime="00:01:23.65" resultid="2317" heatid="6403" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Korona Kraków C 1" number="1">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+77" swimtime="00:01:53.50" resultid="2332" heatid="6533" lane="5" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:00:56.67" />
                    <SPLIT distance="150" swimtime="00:01:24.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2189" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2225" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="2182" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="2255" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Korona Kraków E" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+90" swimtime="00:02:57.42" resultid="2331" heatid="6523" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.72" />
                    <SPLIT distance="100" swimtime="00:01:26.40" />
                    <SPLIT distance="150" swimtime="00:02:13.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2229" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="2244" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2203" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="2196" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Korona Kraków C 1" number="2">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+67" swimtime="00:02:05.91" resultid="2328" heatid="6525" lane="2" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="100" swimtime="00:01:05.42" />
                    <SPLIT distance="150" swimtime="00:01:36.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2189" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="2225" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="2182" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="2255" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Korona Kraków C 2" number="2">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+92" swimtime="00:02:10.40" resultid="2329" heatid="6531" lane="3" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:06.60" />
                    <SPLIT distance="150" swimtime="00:01:39.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2166" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="2269" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2314" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="2185" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Korona Kraków C 2" number="3">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+71" swimtime="00:02:25.91" resultid="2330" heatid="6523" lane="2" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:01:16.06" />
                    <SPLIT distance="150" swimtime="00:01:51.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2185" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="2314" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2166" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2269" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Korona Kraków E" number="3">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+120" swimtime="00:02:27.81" resultid="2333" heatid="6531" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                    <SPLIT distance="150" swimtime="00:01:58.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2196" number="1" reactiontime="+120" />
                    <RELAYPOSITION athleteid="2229" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2203" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2244" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Korona Kraków B" number="1">
              <RESULTS>
                <RESULT eventid="1243" reactiontime="+65" swimtime="00:02:53.23" resultid="2338" heatid="6519" lane="2" entrytime="00:02:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.06" />
                    <SPLIT distance="100" swimtime="00:01:37.64" />
                    <SPLIT distance="150" swimtime="00:02:10.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2259" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2207" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="2276" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="2145" number="4" reactiontime="+86" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Korona Kraków D" number="1">
              <RESULTS>
                <RESULT eventid="1408" reactiontime="+77" swimtime="00:02:17.51" resultid="2334" heatid="6528" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:06.10" />
                    <SPLIT distance="150" swimtime="00:01:41.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2129" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2136" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2141" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="2217" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="Korona Kraków C" number="2">
              <RESULTS>
                <RESULT eventid="1408" reactiontime="+112" swimtime="00:03:06.52" resultid="2335" heatid="6527" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.57" />
                    <SPLIT distance="100" swimtime="00:01:39.04" />
                    <SPLIT distance="150" swimtime="00:02:24.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2259" number="1" reactiontime="+112" />
                    <RELAYPOSITION athleteid="2153" number="2" reactiontime="+110" />
                    <RELAYPOSITION athleteid="2145" number="3" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2193" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1243" reactiontime="+66" swimtime="00:02:21.85" resultid="2336" heatid="6520" lane="4" entrytime="00:02:18.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:15.78" />
                    <SPLIT distance="150" swimtime="00:01:50.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2237" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2141" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="2136" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="2129" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Korona Kraków B" number="3">
              <RESULTS>
                <RESULT eventid="1408" reactiontime="+71" swimtime="00:02:14.31" resultid="2337" heatid="6528" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                    <SPLIT distance="100" swimtime="00:01:08.00" />
                    <SPLIT distance="150" swimtime="00:01:43.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2237" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="2309" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2207" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="2276" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Korona Kraków D" number="3">
              <RESULTS>
                <RESULT eventid="1243" reactiontime="+72" swimtime="00:02:52.87" resultid="2339" heatid="6519" lane="3" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                    <SPLIT distance="100" swimtime="00:01:36.55" />
                    <SPLIT distance="150" swimtime="00:02:16.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2217" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="2153" number="2" reactiontime="+91" />
                    <RELAYPOSITION athleteid="2290" number="3" reactiontime="+93" />
                    <RELAYPOSITION athleteid="2309" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Korona Kraków B" number="1">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+77" swimtime="00:02:04.11" resultid="2318" heatid="6497" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                    <SPLIT distance="100" swimtime="00:01:04.77" />
                    <SPLIT distance="150" swimtime="00:01:39.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2276" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2309" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="2255" number="3" reactiontime="+143" />
                    <RELAYPOSITION athleteid="2307" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Korona Kraków C" number="2">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+75" swimtime="00:01:56.63" resultid="2320" heatid="6497" lane="4" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                    <SPLIT distance="100" swimtime="00:00:56.54" />
                    <SPLIT distance="150" swimtime="00:01:27.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2237" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="2189" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="2129" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2244" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Korona Kraków D 1" number="3">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+89" swimtime="00:02:09.08" resultid="2319" heatid="6496" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:05.07" />
                    <SPLIT distance="150" swimtime="00:01:33.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2141" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="2166" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="2182" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="2217" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Korona Kraków E" number="4">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+108" swimtime="00:02:37.40" resultid="2321" heatid="6495" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.54" />
                    <SPLIT distance="100" swimtime="00:01:20.18" />
                    <SPLIT distance="150" swimtime="00:02:05.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2196" number="1" reactiontime="+108" />
                    <RELAYPOSITION athleteid="2136" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="2153" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="2229" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Korona Kraków  D 2" number="5">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+109" swimtime="00:02:46.07" resultid="2322" heatid="6495" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:36.42" />
                    <SPLIT distance="150" swimtime="00:02:12.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2159" number="1" reactiontime="+109" />
                    <RELAYPOSITION athleteid="2203" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="2207" number="3" />
                    <RELAYPOSITION athleteid="2269" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Korona Kraków B" number="6">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+80" swimtime="00:02:14.17" resultid="2323" heatid="6538" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="100" swimtime="00:01:12.42" />
                    <SPLIT distance="150" swimtime="00:01:42.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2237" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2276" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="2182" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="2266" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Korona Kraków C" number="7">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+62" swimtime="00:02:13.41" resultid="2324" heatid="6538" lane="4" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:11.79" />
                    <SPLIT distance="150" swimtime="00:01:47.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2129" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="2225" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="2136" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="2307" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Korona Kraków D 1" number="8">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+69" swimtime="00:02:19.07" resultid="2325" heatid="6537" lane="2" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                    <SPLIT distance="150" swimtime="00:01:43.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2189" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2141" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="2244" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2217" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Korona Kraków D2" number="9">
              <RESULTS>
                <RESULT eventid="1588" status="DNS" swimtime="00:00:00.00" resultid="2326" heatid="6536" lane="1" entrytime="00:02:45.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2290" number="1" />
                    <RELAYPOSITION athleteid="2159" number="2" />
                    <RELAYPOSITION athleteid="2166" number="3" />
                    <RELAYPOSITION athleteid="2269" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Korona Kraków E" number="10">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+77" swimtime="00:03:11.37" resultid="2327" heatid="6536" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.33" />
                    <SPLIT distance="100" swimtime="00:01:44.68" />
                    <SPLIT distance="150" swimtime="00:02:26.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2309" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2153" number="2" reactiontime="+105" />
                    <RELAYPOSITION athleteid="2229" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2196" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02914" name="UKS Victoria Józefów" nation="POL" region="MAZ">
          <CONTACT email="ali90@o2.pl" name="kowalczyk alicja" />
          <ATHLETES>
            <ATHLETE birthdate="1966-03-01" firstname="Jan" gender="M" lastname="Kośmider" nation="POL" athleteid="2378">
              <RESULTS>
                <RESULT eventid="1092" points="620" reactiontime="+87" swimtime="00:05:56.17" resultid="2379" heatid="6491" lane="5" entrytime="00:05:45.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:05.66" />
                    <SPLIT distance="200" swimtime="00:02:51.00" />
                    <SPLIT distance="250" swimtime="00:03:39.74" />
                    <SPLIT distance="300" swimtime="00:04:30.02" />
                    <SPLIT distance="350" swimtime="00:05:13.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="2380" heatid="6116" lane="6" entrytime="00:02:50.54" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="2381" heatid="6172" lane="3" entrytime="00:01:02.04" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="2382" heatid="6212" lane="3" entrytime="00:00:36.50" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="2383" heatid="6287" lane="2" entrytime="00:02:20.09" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="2384" heatid="6355" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="1610" status="DNS" swimtime="00:00:00.00" resultid="2385" heatid="6405" lane="4" entrytime="00:01:18.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-11-08" firstname="Alicja" gender="F" lastname="Kowalczyk-Kędzierska" nation="POL" athleteid="2386">
              <RESULTS>
                <RESULT eventid="1058" points="472" reactiontime="+88" swimtime="00:06:24.28" resultid="2387" heatid="6430" lane="6" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                    <SPLIT distance="100" swimtime="00:01:31.17" />
                    <SPLIT distance="150" swimtime="00:02:19.28" />
                    <SPLIT distance="200" swimtime="00:03:09.14" />
                    <SPLIT distance="250" swimtime="00:04:03.24" />
                    <SPLIT distance="300" swimtime="00:04:58.23" />
                    <SPLIT distance="350" swimtime="00:05:42.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="470" reactiontime="+89" swimtime="00:01:23.62" resultid="2388" heatid="6080" lane="4" entrytime="00:01:22.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="519" reactiontime="+93" swimtime="00:00:37.92" resultid="2389" heatid="6124" lane="1" entrytime="00:00:37.49" />
                <RESULT eventid="1348" points="559" swimtime="00:00:35.00" resultid="2390" heatid="6221" lane="2" entrytime="00:00:35.20" />
                <RESULT eventid="1378" points="507" reactiontime="+88" swimtime="00:01:22.14" resultid="2391" heatid="6247" lane="2" entrytime="00:01:22.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="405" reactiontime="+90" swimtime="00:01:26.41" resultid="2392" heatid="6314" lane="3" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="484" reactiontime="+93" swimtime="00:02:57.10" resultid="2393" heatid="6370" lane="1" entrytime="00:03:09.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                    <SPLIT distance="100" swimtime="00:01:27.59" />
                    <SPLIT distance="150" swimtime="00:02:13.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Radlin" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1976-01-01" firstname="Dariusz" gender="M" lastname="Krause" nation="POL" athleteid="2395">
              <RESULTS>
                <RESULT eventid="1168" points="306" reactiontime="+82" swimtime="00:01:26.66" resultid="2396" heatid="6087" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="380" reactiontime="+75" swimtime="00:01:10.98" resultid="2397" heatid="6163" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="442" reactiontime="+88" swimtime="00:00:30.39" resultid="2398" heatid="6348" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1640" points="263" reactiontime="+101" swimtime="00:06:22.83" resultid="2399" heatid="6563" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:21.58" />
                    <SPLIT distance="150" swimtime="00:02:09.34" />
                    <SPLIT distance="200" swimtime="00:02:59.11" />
                    <SPLIT distance="250" swimtime="00:03:49.37" />
                    <SPLIT distance="300" swimtime="00:04:41.57" />
                    <SPLIT distance="350" swimtime="00:05:33.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KSWAR" name="KS Warta Poznań" nation="POL" region="WIE">
          <CONTACT city="Poznań" email="j.thiem@glos.com" name="Thiem Jacek" phone="502499565" state="WLKP" street="Os. Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1963-02-17" firstname="JACEK" gender="M" lastname="THIEM" nation="POL" license="MOO11520005" athleteid="2401">
              <RESULTS>
                <RESULT eventid="1092" points="411" reactiontime="+106" swimtime="00:06:48.48" resultid="2402" heatid="6488" lane="2" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:28.32" />
                    <SPLIT distance="150" swimtime="00:02:25.73" />
                    <SPLIT distance="200" swimtime="00:03:21.57" />
                    <SPLIT distance="250" swimtime="00:04:19.95" />
                    <SPLIT distance="300" swimtime="00:05:20.79" />
                    <SPLIT distance="350" swimtime="00:06:06.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="492" reactiontime="+104" swimtime="00:02:59.51" resultid="2403" heatid="6187" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:26.74" />
                    <SPLIT distance="150" swimtime="00:02:12.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="406" reactiontime="+96" swimtime="00:00:36.98" resultid="2404" heatid="6227" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1437" points="450" swimtime="00:02:39.88" resultid="2405" heatid="6282" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:01:19.68" />
                    <SPLIT distance="150" swimtime="00:02:01.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="456" reactiontime="+103" swimtime="00:01:19.67" resultid="2406" heatid="6320" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="425" reactiontime="+108" swimtime="00:05:49.37" resultid="2407" heatid="6564" lane="2" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:25.07" />
                    <SPLIT distance="150" swimtime="00:02:09.72" />
                    <SPLIT distance="200" swimtime="00:02:55.35" />
                    <SPLIT distance="250" swimtime="00:03:40.04" />
                    <SPLIT distance="300" swimtime="00:04:24.37" />
                    <SPLIT distance="350" swimtime="00:05:08.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="ANNA" gender="F" lastname="KOTECKA" nation="POL" athleteid="2408">
              <RESULTS>
                <RESULT eventid="1122" points="513" swimtime="00:12:49.95" resultid="2409" heatid="6444" lane="1" entrytime="00:12:45.00">
                  <SPLITS>
                    <SPLIT distance="400" swimtime="00:06:15.18" />
                    <SPLIT distance="500" swimtime="00:07:54.14" />
                    <SPLIT distance="600" swimtime="00:09:33.36" />
                    <SPLIT distance="700" swimtime="00:11:13.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="393" reactiontime="+90" swimtime="00:00:45.54" resultid="2410" heatid="6121" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="1257" points="492" swimtime="00:01:20.45" resultid="2411" heatid="6153" lane="3" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="445" reactiontime="+89" swimtime="00:01:35.75" resultid="2412" heatid="6246" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="478" swimtime="00:02:56.43" resultid="2413" heatid="6275" lane="4" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                    <SPLIT distance="100" swimtime="00:01:23.65" />
                    <SPLIT distance="150" swimtime="00:02:09.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="539" reactiontime="+91" swimtime="00:03:19.50" resultid="2414" heatid="6369" lane="5" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.20" />
                    <SPLIT distance="100" swimtime="00:01:37.03" />
                    <SPLIT distance="150" swimtime="00:02:29.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="494" swimtime="00:06:10.36" resultid="2415" heatid="6556" lane="4" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:01:25.87" />
                    <SPLIT distance="150" swimtime="00:02:12.18" />
                    <SPLIT distance="200" swimtime="00:02:59.03" />
                    <SPLIT distance="250" swimtime="00:03:46.40" />
                    <SPLIT distance="300" swimtime="00:04:34.70" />
                    <SPLIT distance="350" swimtime="00:05:23.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-17" firstname="REMIGIUSZ" gender="M" lastname="GRZEŚKOWIAK" nation="POL" athleteid="2416">
              <RESULTS>
                <RESULT eventid="1228" points="517" reactiontime="+83" swimtime="00:00:31.69" resultid="2417" heatid="6138" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1272" points="551" reactiontime="+80" swimtime="00:01:00.23" resultid="2418" heatid="6176" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="602" reactiontime="+75" swimtime="00:00:26.42" resultid="2419" heatid="6362" lane="1" entrytime="00:00:26.30" />
                <RESULT eventid="1640" points="458" reactiontime="+76" swimtime="00:05:02.10" resultid="2420" heatid="6570" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:06.84" />
                    <SPLIT distance="150" swimtime="00:01:45.41" />
                    <SPLIT distance="200" swimtime="00:02:24.55" />
                    <SPLIT distance="250" swimtime="00:03:05.65" />
                    <SPLIT distance="300" swimtime="00:03:45.76" />
                    <SPLIT distance="350" swimtime="00:04:25.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-18" firstname="JAKUB" gender="M" lastname="ROMEL" nation="POL" athleteid="2421">
              <RESULTS>
                <RESULT eventid="1092" points="661" reactiontime="+67" swimtime="00:05:12.10" resultid="2422" heatid="6492" lane="5" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:07.91" />
                    <SPLIT distance="150" swimtime="00:01:47.72" />
                    <SPLIT distance="200" swimtime="00:02:27.76" />
                    <SPLIT distance="250" swimtime="00:03:12.68" />
                    <SPLIT distance="300" swimtime="00:03:59.31" />
                    <SPLIT distance="350" swimtime="00:04:36.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="662" reactiontime="+68" swimtime="00:02:24.41" resultid="2423" heatid="6190" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:09.24" />
                    <SPLIT distance="150" swimtime="00:01:46.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="557" reactiontime="+67" swimtime="00:02:14.46" resultid="2424" heatid="6290" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="100" swimtime="00:01:04.48" />
                    <SPLIT distance="150" swimtime="00:01:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" status="DNS" swimtime="00:00:00.00" resultid="2425" heatid="6569" lane="4" entrytime="00:04:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="DARIUSZ" gender="M" lastname="JANYGA" nation="POL" license="M0011520006" athleteid="2426">
              <RESULTS>
                <RESULT eventid="1228" points="619" reactiontime="+92" swimtime="00:00:33.86" resultid="2427" heatid="6132" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1272" points="618" reactiontime="+88" swimtime="00:01:04.29" resultid="2428" heatid="6169" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="698" reactiontime="+54" swimtime="00:01:13.33" resultid="2429" heatid="6258" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="625" reactiontime="+89" swimtime="00:00:28.68" resultid="2430" heatid="6353" lane="4" entrytime="00:00:29.20" />
                <RESULT eventid="1558" points="611" reactiontime="+79" swimtime="00:02:46.01" resultid="2431" heatid="6378" lane="2" entrytime="00:02:50.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:20.91" />
                    <SPLIT distance="150" swimtime="00:02:03.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-02" firstname="PAWEŁ" gender="M" lastname="OLSZEWSKI" nation="POL" license="MOO11520003" athleteid="2432">
              <RESULTS>
                <RESULT eventid="1272" points="843" reactiontime="+76" swimtime="00:01:00.21" resultid="2433" heatid="6173" lane="1" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="775" reactiontime="+76" swimtime="00:02:15.33" resultid="2434" heatid="6288" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="100" swimtime="00:01:05.99" />
                    <SPLIT distance="150" swimtime="00:01:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="799" reactiontime="+76" swimtime="00:00:27.34" resultid="2435" heatid="6356" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1640" points="751" reactiontime="+87" swimtime="00:04:55.24" resultid="2436" heatid="6568" lane="2" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:09.81" />
                    <SPLIT distance="150" swimtime="00:01:46.68" />
                    <SPLIT distance="200" swimtime="00:02:24.72" />
                    <SPLIT distance="250" swimtime="00:03:03.14" />
                    <SPLIT distance="300" swimtime="00:03:41.68" />
                    <SPLIT distance="350" swimtime="00:04:19.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-17" firstname="RADOSŁAW" gender="M" lastname="SOBKOWIAK" nation="POL" athleteid="2437">
              <RESULTS>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="2438" heatid="6162" lane="1" entrytime="00:01:20.00" />
                <RESULT eventid="1528" points="394" reactiontime="+96" swimtime="00:00:31.56" resultid="2439" heatid="6351" lane="5" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="ADRIAN" gender="M" lastname="SOBKOWIAK" nation="POL" athleteid="2440">
              <RESULTS>
                <RESULT eventid="1168" points="379" reactiontime="+99" swimtime="00:01:25.25" resultid="2441" heatid="6088" lane="6" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="341" reactiontime="+88" swimtime="00:00:42.19" resultid="2442" heatid="6209" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1363" status="DNS" swimtime="00:00:00.00" resultid="2443" heatid="6226" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1610" points="366" reactiontime="+88" swimtime="00:01:33.90" resultid="2444" heatid="6399" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="KU AZS UR Kraków" nation="POL">
          <CONTACT city="Kraków" name="Nawrocka" phone="606704926" street="Stańczyka" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-15" firstname="Manuela" gender="F" lastname="Nawrocka" nation="POL" athleteid="2446">
              <RESULTS>
                <RESULT eventid="1153" points="713" reactiontime="+84" swimtime="00:01:14.97" resultid="2447" heatid="6082" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="585" reactiontime="+70" swimtime="00:00:35.60" resultid="2448" heatid="6125" lane="4" entrytime="00:00:33.80" />
                <RESULT eventid="1348" points="496" reactiontime="+82" swimtime="00:00:34.85" resultid="2449" heatid="6222" lane="6" entrytime="00:00:34.60" />
                <RESULT eventid="1452" points="588" reactiontime="+87" swimtime="00:02:45.76" resultid="2450" heatid="6298" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:20.45" />
                    <SPLIT distance="150" swimtime="00:02:08.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="605" reactiontime="+79" swimtime="00:00:30.28" resultid="2451" heatid="6339" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1543" points="557" reactiontime="+72" swimtime="00:02:44.79" resultid="2452" heatid="6371" lane="2" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:19.64" />
                    <SPLIT distance="150" swimtime="00:02:01.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="UKS Wodnik Siemianowice" nation="POL" region="SLA">
          <CONTACT city="Siemianowice Śl." email="mlisienski@all.pl" internet="www.ukswodnik.pl" name="UKS Wodnik Siemianowice" phone="695452707" state="ŚLĄSK" street="Mikołaja 3" zip="41-106" />
          <ATHLETES>
            <ATHLETE birthdate="1987-03-18" firstname="Michał" gender="M" lastname="Lisieński" nation="POL" athleteid="2454">
              <RESULTS>
                <RESULT eventid="1092" points="650" reactiontime="+85" swimtime="00:05:13.75" resultid="2455" heatid="6491" lane="4" entrytime="00:05:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:07.88" />
                    <SPLIT distance="150" swimtime="00:01:48.93" />
                    <SPLIT distance="200" swimtime="00:02:28.78" />
                    <SPLIT distance="250" swimtime="00:03:14.89" />
                    <SPLIT distance="300" swimtime="00:04:00.35" />
                    <SPLIT distance="350" swimtime="00:04:37.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="630" reactiontime="+79" swimtime="00:01:04.77" resultid="2456" heatid="6323" lane="4" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="S02401" name="Miejski Klub Pływacki &quot;ATOL&quot; Oleśnica" nation="POL" region="DOL" shortname="Miejski Klub Pływacki &quot;ATOL&quot; O">
          <CONTACT city="Oleśnica" email="mkp.atol@wp.pl" name="Salik" phone="793018283" state="DOL" street="Przyjaźni" zip="56-400" />
          <ATHLETES>
            <ATHLETE birthdate="1980-02-06" firstname="Marcin" gender="M" lastname="Hejninger" nation="POL" athleteid="2458">
              <RESULTS>
                <RESULT eventid="1333" points="439" reactiontime="+90" swimtime="00:00:38.74" resultid="2459" heatid="6205" lane="4" entrytime="00:00:45.13" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-28" firstname="Marta" gender="F" lastname="Skorek" nation="POL" athleteid="2460">
              <RESULTS>
                <RESULT eventid="1318" points="232" reactiontime="+101" swimtime="00:00:55.43" resultid="2461" heatid="6197" lane="6" entrytime="00:00:49.94" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" name="MOTYL SENIOR MOSiR Stalowa Wola" nation="POL" region="PDK" shortname="MOTYL SENIOR MOSiR Stalowa Wol">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" phone="15-8422562 wew.45" state="PODK." street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1970-06-07" firstname="Wiesław" gender="M" lastname="Bar" nation="POL" athleteid="2473">
              <RESULTS>
                <RESULT eventid="1137" points="505" swimtime="00:10:50.04" resultid="2474" heatid="6454" lane="5" entrytime="00:11:01.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:10.17" />
                    <SPLIT distance="200" swimtime="00:02:28.18" />
                    <SPLIT distance="300" swimtime="00:03:48.68" />
                    <SPLIT distance="400" swimtime="00:05:10.93" />
                    <SPLIT distance="500" swimtime="00:06:33.96" />
                    <SPLIT distance="600" swimtime="00:07:59.40" />
                    <SPLIT distance="700" swimtime="00:09:24.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="621" reactiontime="+90" swimtime="00:01:12.35" resultid="2475" heatid="6093" lane="2" entrytime="00:01:13.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - przedwczesny start" eventid="1272" reactiontime="+75" status="DSQ" swimtime="00:01:01.64" resultid="2476" heatid="6173" lane="5" entrytime="00:01:01.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="579" reactiontime="+91" swimtime="00:02:21.99" resultid="2477" heatid="6288" lane="1" entrytime="00:02:18.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:09.54" />
                    <SPLIT distance="150" swimtime="00:01:45.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="595" reactiontime="+90" swimtime="00:02:42.11" resultid="2478" heatid="6307" lane="3" entrytime="00:02:41.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:16.69" />
                    <SPLIT distance="150" swimtime="00:02:06.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="692" reactiontime="+81" swimtime="00:00:27.60" resultid="2479" heatid="6359" lane="5" entrytime="00:00:27.44" />
                <RESULT eventid="1640" points="554" reactiontime="+92" swimtime="00:05:05.84" resultid="2480" heatid="6567" lane="1" entrytime="00:05:03.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                    <SPLIT distance="150" swimtime="00:01:47.48" />
                    <SPLIT distance="200" swimtime="00:02:26.17" />
                    <SPLIT distance="250" swimtime="00:03:05.62" />
                    <SPLIT distance="300" swimtime="00:03:45.60" />
                    <SPLIT distance="350" swimtime="00:04:26.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="Baran" nation="POL" athleteid="2481">
              <RESULTS>
                <RESULT eventid="1228" points="759" reactiontime="+77" swimtime="00:00:30.12" resultid="2482" heatid="6138" lane="3" entrytime="00:00:29.94" />
                <RESULT eventid="1272" points="651" reactiontime="+87" swimtime="00:00:59.34" resultid="2483" heatid="6177" lane="6" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="507" reactiontime="+88" swimtime="00:00:31.52" resultid="2484" heatid="6234" lane="3" entrytime="00:00:30.66" />
                <RESULT eventid="1393" points="722" reactiontime="+75" swimtime="00:01:05.54" resultid="2485" heatid="6261" lane="3" entrytime="00:01:05.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="652" reactiontime="+75" swimtime="00:00:26.69" resultid="2486" heatid="6361" lane="3" entrytime="00:00:26.50" />
                <RESULT eventid="1558" points="633" reactiontime="+74" swimtime="00:02:28.06" resultid="2487" heatid="6381" lane="4" entrytime="00:02:25.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="2488">
              <RESULTS>
                <RESULT eventid="1092" points="824" reactiontime="+75" swimtime="00:05:04.39" resultid="2489" heatid="6492" lane="3" entrytime="00:05:05.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:06.91" />
                    <SPLIT distance="150" swimtime="00:01:46.40" />
                    <SPLIT distance="200" swimtime="00:02:25.25" />
                    <SPLIT distance="250" swimtime="00:03:08.12" />
                    <SPLIT distance="300" swimtime="00:03:51.13" />
                    <SPLIT distance="350" swimtime="00:04:28.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="725" reactiontime="+77" swimtime="00:01:05.00" resultid="2490" heatid="6099" lane="1" entrytime="00:01:04.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="773" reactiontime="+77" swimtime="00:02:21.46" resultid="2491" heatid="6191" lane="5" entrytime="00:02:20.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="771" reactiontime="+74" swimtime="00:02:06.67" resultid="2492" heatid="6292" lane="6" entrytime="00:02:04.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                    <SPLIT distance="100" swimtime="00:01:00.07" />
                    <SPLIT distance="150" swimtime="00:01:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="681" reactiontime="+75" swimtime="00:02:22.51" resultid="2493" heatid="6311" lane="1" entrytime="00:02:20.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:07.07" />
                    <SPLIT distance="150" swimtime="00:01:48.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="852" reactiontime="+73" swimtime="00:01:00.20" resultid="2494" heatid="6326" lane="3" entrytime="00:01:00.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="735" reactiontime="+76" swimtime="00:04:31.86" resultid="2495" heatid="6570" lane="1" entrytime="00:04:29.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                    <SPLIT distance="100" swimtime="00:01:03.38" />
                    <SPLIT distance="150" swimtime="00:01:37.42" />
                    <SPLIT distance="200" swimtime="00:02:12.20" />
                    <SPLIT distance="250" swimtime="00:02:47.12" />
                    <SPLIT distance="300" swimtime="00:03:22.11" />
                    <SPLIT distance="350" swimtime="00:03:57.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Paweł" gender="M" lastname="Cieśliński" nation="POL" athleteid="2496">
              <RESULTS>
                <RESULT eventid="1137" points="298" swimtime="00:12:50.35" resultid="2497" heatid="6450" lane="5" entrytime="00:12:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:26.74" />
                    <SPLIT distance="200" swimtime="00:03:00.65" />
                    <SPLIT distance="300" swimtime="00:04:40.33" />
                    <SPLIT distance="400" swimtime="00:06:19.42" />
                    <SPLIT distance="500" swimtime="00:07:57.52" />
                    <SPLIT distance="600" swimtime="00:09:36.53" />
                    <SPLIT distance="700" swimtime="00:11:14.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="493" reactiontime="+89" swimtime="00:02:59.49" resultid="2498" heatid="6113" lane="2" entrytime="00:03:05.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:01:26.41" />
                    <SPLIT distance="150" swimtime="00:02:13.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="355" reactiontime="+103" swimtime="00:03:03.36" resultid="2499" heatid="6188" lane="6" entrytime="00:03:05.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:27.93" />
                    <SPLIT distance="150" swimtime="00:02:16.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="442" reactiontime="+83" swimtime="00:00:37.80" resultid="2500" heatid="6212" lane="5" entrytime="00:00:37.01" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="2501" heatid="6304" lane="3" entrytime="00:02:57.00" />
                <RESULT eventid="1610" points="430" reactiontime="+87" swimtime="00:01:23.80" resultid="2502" heatid="6404" lane="5" entrytime="00:01:21.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-07" firstname="Paweł" gender="M" lastname="Ciurko" nation="POL" athleteid="2503">
              <RESULTS>
                <RESULT eventid="1092" points="386" reactiontime="+93" swimtime="00:06:17.03" resultid="2504" heatid="6490" lane="3" entrytime="00:06:01.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:01:27.70" />
                    <SPLIT distance="150" swimtime="00:02:21.13" />
                    <SPLIT distance="200" swimtime="00:03:14.64" />
                    <SPLIT distance="250" swimtime="00:04:01.59" />
                    <SPLIT distance="300" swimtime="00:04:50.59" />
                    <SPLIT distance="350" swimtime="00:05:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="516" reactiontime="+92" swimtime="00:02:55.17" resultid="2505" heatid="6116" lane="1" entrytime="00:02:48.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.60" />
                    <SPLIT distance="100" swimtime="00:01:22.17" />
                    <SPLIT distance="150" swimtime="00:02:08.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="283" reactiontime="+95" swimtime="00:03:11.51" resultid="2506" heatid="6189" lane="5" entrytime="00:02:58.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                    <SPLIT distance="100" swimtime="00:01:31.64" />
                    <SPLIT distance="150" swimtime="00:02:21.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="287" reactiontime="+91" swimtime="00:00:38.28" resultid="2507" heatid="6230" lane="4" entrytime="00:00:33.02" />
                <RESULT eventid="1467" points="423" reactiontime="+89" swimtime="00:02:51.39" resultid="2508" heatid="6307" lane="1" entrytime="00:02:47.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:25.63" />
                    <SPLIT distance="150" swimtime="00:02:11.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="364" reactiontime="+87" swimtime="00:01:17.97" resultid="2509" heatid="6321" lane="5" entrytime="00:01:19.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="552" reactiontime="+89" swimtime="00:01:19.07" resultid="2510" heatid="6406" lane="3" entrytime="00:01:15.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-09" firstname="Włodzimierz" gender="M" lastname="Jarzyna" nation="POL" athleteid="2511">
              <RESULTS>
                <RESULT eventid="1092" points="570" reactiontime="+96" swimtime="00:06:59.95" resultid="2512" heatid="6487" lane="5" entrytime="00:07:25.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                    <SPLIT distance="100" swimtime="00:01:44.54" />
                    <SPLIT distance="150" swimtime="00:03:31.07" />
                    <SPLIT distance="200" swimtime="00:04:30.36" />
                    <SPLIT distance="250" swimtime="00:05:29.64" />
                    <SPLIT distance="300" swimtime="00:06:16.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="562" reactiontime="+97" swimtime="00:01:27.10" resultid="2513" heatid="6086" lane="6" entrytime="00:01:36.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="559" reactiontime="+91" swimtime="00:03:34.27" resultid="2514" heatid="6110" lane="4" entrytime="00:03:41.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="100" swimtime="00:01:43.97" />
                    <SPLIT distance="150" swimtime="00:02:41.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="547" reactiontime="+72" swimtime="00:01:29.97" resultid="2515" heatid="6253" lane="6" entrytime="00:01:36.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="519" reactiontime="+96" swimtime="00:03:20.48" resultid="2516" heatid="6301" lane="4" entrytime="00:03:38.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                    <SPLIT distance="100" swimtime="00:01:36.06" />
                    <SPLIT distance="150" swimtime="00:02:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="527" reactiontime="+78" swimtime="00:03:20.34" resultid="2517" heatid="6374" lane="3" entrytime="00:03:36.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                    <SPLIT distance="100" swimtime="00:01:39.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="474" reactiontime="+101" swimtime="00:06:18.37" resultid="2518" heatid="6562" lane="5" entrytime="00:06:24.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:30.02" />
                    <SPLIT distance="150" swimtime="00:02:19.43" />
                    <SPLIT distance="200" swimtime="00:03:09.44" />
                    <SPLIT distance="250" swimtime="00:03:58.09" />
                    <SPLIT distance="300" swimtime="00:04:46.66" />
                    <SPLIT distance="350" swimtime="00:05:34.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-18" firstname="Waldemar" gender="M" lastname="Kalbarczyk" nation="POL" athleteid="2519">
              <RESULTS>
                <RESULT eventid="1092" points="495" reactiontime="+87" swimtime="00:06:10.81" resultid="2520" heatid="6489" lane="2" entrytime="00:06:18.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:22.44" />
                    <SPLIT distance="150" swimtime="00:02:08.50" />
                    <SPLIT distance="200" swimtime="00:02:54.30" />
                    <SPLIT distance="250" swimtime="00:03:46.70" />
                    <SPLIT distance="300" swimtime="00:04:40.91" />
                    <SPLIT distance="350" swimtime="00:05:25.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="536" reactiontime="+85" swimtime="00:01:15.98" resultid="2521" heatid="6092" lane="6" entrytime="00:01:16.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="479" reactiontime="+89" swimtime="00:01:08.25" resultid="2522" heatid="6170" lane="5" entrytime="00:01:05.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="465" reactiontime="+68" swimtime="00:01:18.37" resultid="2523" heatid="6256" lane="6" entrytime="00:01:21.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="512" reactiontime="+83" swimtime="00:02:50.37" resultid="2524" heatid="6305" lane="3" entrytime="00:02:51.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:20.52" />
                    <SPLIT distance="150" swimtime="00:02:10.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="579" reactiontime="+82" swimtime="00:00:29.29" resultid="2525" heatid="6353" lane="2" entrytime="00:00:29.31" />
                <RESULT eventid="1558" points="506" reactiontime="+79" swimtime="00:02:49.98" resultid="2526" heatid="6377" lane="2" entrytime="00:02:55.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:24.10" />
                    <SPLIT distance="150" swimtime="00:02:08.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="2527">
              <RESULTS>
                <RESULT eventid="1092" points="636" reactiontime="+87" swimtime="00:06:07.70" resultid="2528" heatid="6489" lane="4" entrytime="00:06:13.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="100" swimtime="00:01:23.18" />
                    <SPLIT distance="150" swimtime="00:02:09.30" />
                    <SPLIT distance="200" swimtime="00:02:55.70" />
                    <SPLIT distance="250" swimtime="00:03:50.65" />
                    <SPLIT distance="300" swimtime="00:04:44.59" />
                    <SPLIT distance="350" swimtime="00:05:27.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="586" reactiontime="+87" swimtime="00:01:07.98" resultid="2529" heatid="6168" lane="4" entrytime="00:01:08.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="481" reactiontime="+92" swimtime="00:03:11.69" resultid="2530" heatid="6187" lane="2" entrytime="00:03:10.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:30.72" />
                    <SPLIT distance="150" swimtime="00:02:23.49" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - przedwczesny start." eventid="1437" reactiontime="+41" status="DSQ" swimtime="00:02:33.81" resultid="2531" heatid="6285" lane="5" entrytime="00:02:32.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:12.65" />
                    <SPLIT distance="150" swimtime="00:01:53.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="606" reactiontime="+91" swimtime="00:02:55.52" resultid="2532" heatid="6306" lane="6" entrytime="00:02:51.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:23.78" />
                    <SPLIT distance="150" swimtime="00:02:17.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="492" reactiontime="+84" swimtime="00:01:20.01" resultid="2533" heatid="6320" lane="2" entrytime="00:01:22.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="594" reactiontime="+87" swimtime="00:02:57.17" resultid="2534" heatid="6377" lane="5" entrytime="00:02:56.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:01:25.52" />
                    <SPLIT distance="150" swimtime="00:02:11.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-11-29" firstname="Jarosław" gender="M" lastname="Niedbałowski" nation="POL" athleteid="2535">
              <RESULTS>
                <RESULT eventid="1198" points="605" reactiontime="+92" swimtime="00:03:10.56" resultid="2536" heatid="6112" lane="2" entrytime="00:03:15.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:01:28.72" />
                    <SPLIT distance="150" swimtime="00:02:19.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="2537" heatid="6163" lane="3" entrytime="00:01:14.04" />
                <RESULT eventid="1333" points="677" reactiontime="+90" swimtime="00:00:36.66" resultid="2538" heatid="6212" lane="1" entrytime="00:00:37.48" />
                <RESULT eventid="1528" points="505" reactiontime="+81" swimtime="00:00:31.85" resultid="2539" heatid="6350" lane="6" entrytime="00:00:31.42" />
                <RESULT eventid="1610" points="656" reactiontime="+84" swimtime="00:01:23.75" resultid="2540" heatid="6402" lane="2" entrytime="00:01:25.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-04" firstname="Paweł" gender="M" lastname="Opaliński" nation="POL" athleteid="2541">
              <RESULTS>
                <RESULT eventid="1137" points="537" swimtime="00:10:33.62" resultid="2542" heatid="6451" lane="2" entrytime="00:12:00.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:09.80" />
                    <SPLIT distance="200" swimtime="00:02:24.75" />
                    <SPLIT distance="300" swimtime="00:03:43.00" />
                    <SPLIT distance="400" swimtime="00:05:03.21" />
                    <SPLIT distance="500" swimtime="00:06:25.18" />
                    <SPLIT distance="600" swimtime="00:07:47.01" />
                    <SPLIT distance="700" swimtime="00:09:11.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="640" reactiontime="+80" swimtime="00:02:44.48" resultid="2543" heatid="6115" lane="6" entrytime="00:02:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                    <SPLIT distance="150" swimtime="00:02:00.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="631" reactiontime="+83" swimtime="00:00:59.96" resultid="2544" heatid="6174" lane="1" entrytime="00:01:00.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="607" reactiontime="+42" swimtime="00:00:34.02" resultid="2545" heatid="6215" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1437" points="667" reactiontime="+89" swimtime="00:02:12.96" resultid="2546" heatid="6289" lane="4" entrytime="00:02:13.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="590" reactiontime="+80" swimtime="00:01:15.42" resultid="2547" heatid="6407" lane="1" entrytime="00:01:14.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" status="DNS" swimtime="00:00:00.00" resultid="2548" heatid="6567" lane="4" entrytime="00:04:57.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="2549">
              <RESULTS>
                <RESULT eventid="1092" points="477" reactiontime="+81" swimtime="00:06:05.17" resultid="2550" heatid="6490" lane="5" entrytime="00:06:09.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                    <SPLIT distance="100" swimtime="00:01:25.83" />
                    <SPLIT distance="150" swimtime="00:02:13.43" />
                    <SPLIT distance="200" swimtime="00:03:01.44" />
                    <SPLIT distance="250" swimtime="00:03:50.42" />
                    <SPLIT distance="300" swimtime="00:04:40.89" />
                    <SPLIT distance="350" swimtime="00:05:23.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="468" reactiontime="+78" swimtime="00:01:15.17" resultid="2551" heatid="6093" lane="5" entrytime="00:01:13.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="345" reactiontime="+87" swimtime="00:03:05.08" resultid="2552" heatid="6187" lane="6" entrytime="00:03:12.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:29.97" />
                    <SPLIT distance="150" swimtime="00:02:17.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="445" reactiontime="+72" swimtime="00:01:16.99" resultid="2553" heatid="6257" lane="5" entrytime="00:01:16.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="415" reactiontime="+82" swimtime="00:02:48.14" resultid="2554" heatid="6306" lane="3" entrytime="00:02:48.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                    <SPLIT distance="150" swimtime="00:02:09.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="406" reactiontime="+70" swimtime="00:02:51.68" resultid="2555" heatid="6378" lane="5" entrytime="00:02:50.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.72" />
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                    <SPLIT distance="150" swimtime="00:02:10.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="421" reactiontime="+91" swimtime="00:05:27.46" resultid="2556" heatid="6566" lane="6" entrytime="00:05:27.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:16.15" />
                    <SPLIT distance="150" swimtime="00:01:57.74" />
                    <SPLIT distance="200" swimtime="00:02:40.46" />
                    <SPLIT distance="250" swimtime="00:03:23.68" />
                    <SPLIT distance="300" swimtime="00:04:05.99" />
                    <SPLIT distance="350" swimtime="00:04:47.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="2557">
              <RESULTS>
                <RESULT eventid="1058" points="619" reactiontime="+84" swimtime="00:06:43.08" resultid="2558" heatid="6430" lane="3" entrytime="00:06:59.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:01:29.68" />
                    <SPLIT distance="150" swimtime="00:03:17.95" />
                    <SPLIT distance="200" swimtime="00:04:12.73" />
                    <SPLIT distance="250" swimtime="00:05:08.67" />
                    <SPLIT distance="300" swimtime="00:05:56.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="584" reactiontime="+93" swimtime="00:03:24.73" resultid="2559" heatid="6105" lane="3" entrytime="00:03:28.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.58" />
                    <SPLIT distance="100" swimtime="00:01:38.51" />
                    <SPLIT distance="150" swimtime="00:02:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" status="DNS" swimtime="00:00:00.00" resultid="2560" heatid="6154" lane="6" entrytime="00:01:18.02" />
                <RESULT eventid="1348" points="527" reactiontime="+89" swimtime="00:00:37.76" resultid="2561" heatid="6221" lane="6" entrytime="00:00:38.11" />
                <RESULT eventid="1452" points="630" reactiontime="+94" swimtime="00:03:05.51" resultid="2562" heatid="6296" lane="5" entrytime="00:03:11.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:01:32.08" />
                    <SPLIT distance="150" swimtime="00:02:25.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="484" reactiontime="+93" swimtime="00:01:29.57" resultid="2563" heatid="6314" lane="1" entrytime="00:01:35.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="552" reactiontime="+91" swimtime="00:00:34.31" resultid="2564" heatid="6335" lane="2" entrytime="00:00:35.41" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-12" firstname="Adam" gender="M" lastname="Przybylski" nation="POL" athleteid="2565">
              <RESULTS>
                <RESULT eventid="1092" points="479" reactiontime="+90" swimtime="00:06:28.16" resultid="2566" heatid="6489" lane="1" entrytime="00:06:20.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:25.15" />
                    <SPLIT distance="150" swimtime="00:02:14.78" />
                    <SPLIT distance="200" swimtime="00:03:02.91" />
                    <SPLIT distance="250" swimtime="00:04:00.72" />
                    <SPLIT distance="300" swimtime="00:04:58.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="2567" heatid="6133" lane="1" entrytime="00:00:36.12" />
                <RESULT eventid="1302" points="435" reactiontime="+100" swimtime="00:03:07.05" resultid="2568" heatid="6187" lane="5" entrytime="00:03:10.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:01:29.05" />
                    <SPLIT distance="150" swimtime="00:02:18.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="677" reactiontime="+95" swimtime="00:00:31.19" resultid="2569" heatid="6231" lane="3" entrytime="00:00:32.45" />
                <RESULT eventid="1393" points="568" reactiontime="+67" swimtime="00:01:18.55" resultid="2570" heatid="6256" lane="4" entrytime="00:01:18.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="503" reactiontime="+90" swimtime="00:01:17.12" resultid="2571" heatid="6321" lane="2" entrytime="00:01:18.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="533" reactiontime="+68" swimtime="00:02:53.79" resultid="2572" heatid="6377" lane="1" entrytime="00:02:58.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.87" />
                    <SPLIT distance="100" swimtime="00:02:10.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-15" firstname="Michał" gender="M" lastname="Skrok" nation="POL" athleteid="2573">
              <RESULTS>
                <RESULT eventid="1092" points="728" reactiontime="+89" swimtime="00:05:17.25" resultid="2574" heatid="6489" lane="3" entrytime="00:06:10.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:13.06" />
                    <SPLIT distance="150" swimtime="00:01:55.37" />
                    <SPLIT distance="200" swimtime="00:02:36.80" />
                    <SPLIT distance="250" swimtime="00:03:19.54" />
                    <SPLIT distance="300" swimtime="00:04:02.83" />
                    <SPLIT distance="350" swimtime="00:04:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="691" reactiontime="+78" swimtime="00:01:06.03" resultid="2575" heatid="6096" lane="4" entrytime="00:01:08.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. C" eventid="1198" points="721" reactiontime="+76" swimtime="00:02:38.08" resultid="2576" heatid="6115" lane="4" entrytime="00:02:52.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                    <SPLIT distance="150" swimtime="00:01:57.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="697" reactiontime="+76" swimtime="00:00:32.48" resultid="2577" heatid="6215" lane="1" entrytime="00:00:33.70" />
                <RESULT eventid="1467" points="648" reactiontime="+80" swimtime="00:02:24.89" resultid="2578" heatid="6309" lane="3" entrytime="00:02:34.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="150" swimtime="00:01:51.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2579" heatid="6322" lane="3" entrytime="00:01:14.01" />
                <RESULT eventid="1610" points="683" reactiontime="+76" swimtime="00:01:11.85" resultid="2580" heatid="6407" lane="5" entrytime="00:01:14.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-04" firstname="Sebastian" gender="M" lastname="Żarów" nation="POL" athleteid="2581">
              <RESULTS>
                <RESULT eventid="1168" points="442" reactiontime="+84" swimtime="00:01:16.02" resultid="2582" heatid="6090" lane="6" entrytime="00:01:20.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="493" reactiontime="+86" swimtime="00:01:04.00" resultid="2583" heatid="6169" lane="6" entrytime="00:01:07.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="367" reactiontime="+82" swimtime="00:00:39.49" resultid="2584" heatid="6206" lane="4" entrytime="00:00:44.11" />
                <RESULT eventid="1437" points="377" reactiontime="+96" swimtime="00:02:33.11" resultid="2585" heatid="6281" lane="3" entrytime="00:02:45.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:11.06" />
                    <SPLIT distance="150" swimtime="00:01:51.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="487" reactiontime="+86" swimtime="00:00:28.90" resultid="2586" heatid="6353" lane="5" entrytime="00:00:29.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" swimtime="00:01:58.44" resultid="2587" heatid="6526" lane="6" entrytime="00:02:01.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:03.49" />
                    <SPLIT distance="150" swimtime="00:01:31.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2481" number="1" />
                    <RELAYPOSITION athleteid="2573" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="2488" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="2541" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+71" swimtime="00:02:10.85" resultid="2588" heatid="6524" lane="5" entrytime="00:02:15.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:01:43.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2473" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="2503" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="2519" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="2565" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+77" swimtime="00:02:19.57" resultid="2589" heatid="6523" lane="4" entrytime="00:02:22.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:13.86" />
                    <SPLIT distance="150" swimtime="00:01:47.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2527" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2535" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="2549" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="2511" number="4" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+87" swimtime="00:01:50.82" resultid="2590" heatid="6534" lane="1" entrytime="00:01:48.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.23" />
                    <SPLIT distance="100" swimtime="00:00:55.23" />
                    <SPLIT distance="150" swimtime="00:01:22.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2481" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="2573" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="2541" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="2488" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+85" swimtime="00:01:56.55" resultid="2591" heatid="6533" lane="6" entrytime="00:01:56.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="100" swimtime="00:01:01.36" />
                    <SPLIT distance="150" swimtime="00:01:28.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2519" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="2496" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2565" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="2473" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+83" swimtime="00:02:04.27" resultid="2592" heatid="6532" lane="2" entrytime="00:02:02.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="100" swimtime="00:01:02.66" />
                    <SPLIT distance="150" swimtime="00:01:31.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2527" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2535" number="2" />
                    <RELAYPOSITION athleteid="2549" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="2511" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KRK" name="Piotr Urbańczyk" nation="POL" region="MAL">
          <CONTACT city="Kraków" email="piotr_urbanczyk@onet.pl" name="Urbańczyk" phone="608172201" state="MAŁOP" street="os Piastów 57/46" zip="31-625" />
          <ATHLETES>
            <ATHLETE birthdate="1984-03-16" firstname="Piotr" gender="M" lastname="Urbańczyk" nation="POL" athleteid="2628">
              <RESULTS>
                <RESULT eventid="1228" points="712" reactiontime="+76" swimtime="00:00:29.28" resultid="2629" heatid="6139" lane="1" entrytime="00:00:29.07" entrycourse="SCM" />
                <RESULT eventid="1393" points="741" reactiontime="+72" swimtime="00:01:02.12" resultid="2630" heatid="6262" lane="2" entrytime="00:01:00.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="784" reactiontime="+67" swimtime="00:02:15.48" resultid="2631" heatid="6382" lane="4" entrytime="00:02:13.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:06.20" />
                    <SPLIT distance="150" swimtime="00:01:40.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="MOSiR KSZO Ostrowiec Św." nation="POL">
          <CONTACT name="Różalski Józef" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" athleteid="2633">
              <RESULTS>
                <RESULT eventid="1092" points="605" reactiontime="+93" swimtime="00:07:22.03" resultid="2634" heatid="6487" lane="1" entrytime="00:07:30.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                    <SPLIT distance="100" swimtime="00:01:40.80" />
                    <SPLIT distance="150" swimtime="00:02:41.25" />
                    <SPLIT distance="200" swimtime="00:03:41.54" />
                    <SPLIT distance="250" swimtime="00:04:41.52" />
                    <SPLIT distance="300" swimtime="00:05:43.77" />
                    <SPLIT distance="350" swimtime="00:06:33.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="737" reactiontime="+91" swimtime="00:01:23.63" resultid="2635" heatid="6089" lane="2" entrytime="00:01:23.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="744" reactiontime="+89" swimtime="00:01:12.88" resultid="2636" heatid="6165" lane="6" entrytime="00:01:12.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="715" swimtime="00:00:35.61" resultid="2637" heatid="6230" lane="2" entrytime="00:00:33.20" />
                <RESULT eventid="1467" points="583" reactiontime="+96" swimtime="00:03:26.93" resultid="2638" heatid="6302" lane="4" entrytime="00:03:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:39.72" />
                    <SPLIT distance="150" swimtime="00:02:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="535" reactiontime="+96" swimtime="00:01:33.73" resultid="2639" heatid="6319" lane="1" entrytime="00:01:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="724" reactiontime="+90" swimtime="00:00:31.48" resultid="2640" heatid="6350" lane="2" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00305" name="UKS NAWA Skierniewice" nation="POL" region="LOD">
          <CONTACT city="Skierniewice" email="uks_nawa@interia.pl" name="Marcin Sarna" phone="603331973" zip="96-100" />
          <ATHLETES>
            <ATHLETE birthdate="1989-07-11" firstname="Sebastian" gender="M" lastname="Krawczyk" nation="POL" license="S00305200017" athleteid="2642">
              <RESULTS>
                <RESULT eventid="1333" points="821" reactiontime="+84" swimtime="00:00:30.25" resultid="2643" heatid="6217" lane="3" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SMT" name="Szczecin Masters Team" nation="POL" region="ZACHPOM">
          <CONTACT city="szczecin" email="trotyl11@windowslive.com" name="Michal Zaremba" phone="668353622" state="ZACHP" street="Lucznicza 36a/2" zip="71-472" />
          <ATHLETES>
            <ATHLETE birthdate="1988-01-02" firstname="Kamila" gender="F" lastname="Wojdak" nation="POL" athleteid="2645">
              <RESULTS>
                <RESULT eventid="1153" status="DNS" swimtime="00:00:00.00" resultid="2646" heatid="6082" lane="5" entrytime="00:01:14.00" />
                <RESULT eventid="1257" points="671" reactiontime="+86" swimtime="00:01:03.75" resultid="2647" heatid="6158" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="718" reactiontime="+82" swimtime="00:00:36.63" resultid="2648" heatid="6201" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1513" points="661" reactiontime="+84" swimtime="00:00:29.39" resultid="2649" heatid="6340" lane="2" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-22" firstname="Jan" gender="M" lastname="Roening" nation="POL" athleteid="2650">
              <RESULTS>
                <RESULT eventid="1168" points="635" reactiontime="+73" swimtime="00:01:07.37" resultid="2651" heatid="6098" lane="2" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="634" reactiontime="+80" swimtime="00:00:32.93" resultid="2652" heatid="6217" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="1610" points="618" reactiontime="+86" swimtime="00:01:14.15" resultid="2653" heatid="6408" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-22" firstname="Rafal" gender="M" lastname="Lisiecki" nation="POL" athleteid="2654">
              <RESULTS>
                <RESULT eventid="1228" points="548" reactiontime="+73" swimtime="00:00:31.09" resultid="2655" heatid="6137" lane="3" entrytime="00:00:30.30" />
                <RESULT eventid="1393" status="DNS" swimtime="00:00:00.00" resultid="2656" heatid="6259" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1528" points="529" reactiontime="+87" swimtime="00:00:27.59" resultid="2657" heatid="6360" lane="1" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-22" firstname="Szymon" gender="M" lastname="Kluczyk" nation="POL" athleteid="2658">
              <RESULTS>
                <RESULT eventid="1467" points="650" reactiontime="+88" swimtime="00:02:29.02" resultid="2659" heatid="6308" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:54.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-22" firstname="Michal" gender="M" lastname="Zaremba" nation="POL" athleteid="2661">
              <RESULTS>
                <RESULT eventid="1168" points="542" reactiontime="+75" swimtime="00:01:10.99" resultid="2662" heatid="6098" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="549" reactiontime="+80" swimtime="00:02:37.64" resultid="2663" heatid="6309" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:13.99" />
                    <SPLIT distance="150" swimtime="00:02:01.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="523" reactiontime="+78" swimtime="00:01:08.93" resultid="2664" heatid="6324" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-22" firstname="Piotr" gender="M" lastname="Zaremba" nation="POL" athleteid="2665">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="2666" heatid="6099" lane="5" entrytime="00:01:04.00" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="2667" heatid="6310" lane="1" entrytime="00:02:30.00" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2668" heatid="6326" lane="5" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+74" swimtime="00:02:01.27" resultid="2669" heatid="6526" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:03.68" />
                    <SPLIT distance="150" swimtime="00:01:33.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2658" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2661" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2665" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="2650" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Victory Masters Elbląg" nation="POL" region="WAR">
          <CONTACT name="Latecki" />
          <ATHLETES>
            <ATHLETE birthdate="1966-06-06" firstname="Andrzej" gender="M" lastname="Pasieczny" nation="POL" athleteid="2674">
              <RESULTS>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="2675" heatid="6191" lane="1" entrytime="00:02:21.95" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="2676" heatid="6290" lane="5" entrytime="00:02:11.00" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2677" heatid="6325" lane="4" entrytime="00:01:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-12" firstname="Grzegorz" gender="M" lastname="Latecki" nation="POL" athleteid="2679">
              <RESULTS>
                <RESULT eventid="1092" points="725" reactiontime="+81" swimtime="00:05:38.02" resultid="2680" heatid="6491" lane="2" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:16.39" />
                    <SPLIT distance="150" swimtime="00:02:00.48" />
                    <SPLIT distance="200" swimtime="00:02:44.62" />
                    <SPLIT distance="250" swimtime="00:03:32.41" />
                    <SPLIT distance="300" swimtime="00:04:20.91" />
                    <SPLIT distance="350" swimtime="00:05:00.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="710" reactiontime="+69" swimtime="00:00:32.35" resultid="2681" heatid="6136" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1272" points="708" reactiontime="+81" swimtime="00:01:01.44" resultid="2682" heatid="6174" lane="4" entrytime="00:01:00.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="784" reactiontime="+77" swimtime="00:00:29.70" resultid="2683" heatid="6238" lane="6" entrytime="00:00:29.30" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="2684" heatid="6310" lane="6" entrytime="00:02:33.00" />
                <RESULT eventid="1528" points="749" reactiontime="+76" swimtime="00:00:27.00" resultid="2685" heatid="6359" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1558" points="663" reactiontime="+70" swimtime="00:02:41.56" resultid="2686" heatid="6379" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:20.28" />
                    <SPLIT distance="150" swimtime="00:02:02.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-30" firstname="Henryk" gender="M" lastname="Iszoro" nation="POL" athleteid="2687">
              <RESULTS>
                <RESULT eventid="1198" points="331" reactiontime="+116" swimtime="00:04:26.67" resultid="2688" heatid="6109" lane="5" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.62" />
                    <SPLIT distance="100" swimtime="00:02:09.23" />
                    <SPLIT distance="150" swimtime="00:03:20.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="446" reactiontime="+113" swimtime="00:00:47.35" resultid="2689" heatid="6205" lane="1" entrytime="00:00:47.00" />
                <RESULT eventid="1610" points="382" reactiontime="+115" swimtime="00:01:52.15" resultid="2690" heatid="6396" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-09-12" firstname="Tomasz" gender="M" lastname="Gleb" nation="POL" athleteid="2691">
              <RESULTS>
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="2692" heatid="6454" lane="6" entrytime="00:11:15.30" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="2693" heatid="6112" lane="1" entrytime="00:03:20.15" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="2694" heatid="6169" lane="3" entrytime="00:01:06.05" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="2695" heatid="6286" lane="4" entrytime="00:02:25.31" />
                <RESULT eventid="1640" status="DNS" swimtime="00:00:00.00" resultid="2696" heatid="6566" lane="3" entrytime="00:05:15.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="2697">
              <RESULTS>
                <RESULT eventid="1122" points="223" swimtime="00:15:15.70" resultid="2698" heatid="6442" lane="1" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.84" />
                    <SPLIT distance="100" swimtime="00:01:51.20" />
                    <SPLIT distance="200" swimtime="00:03:47.95" />
                    <SPLIT distance="300" swimtime="00:05:44.80" />
                    <SPLIT distance="400" swimtime="00:07:40.60" />
                    <SPLIT distance="500" swimtime="00:09:35.40" />
                    <SPLIT distance="600" swimtime="00:11:29.60" />
                    <SPLIT distance="700" swimtime="00:13:25.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="191" reactiontime="+101" swimtime="00:01:39.66" resultid="2699" heatid="6150" lane="2" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="184" reactiontime="+113" swimtime="00:03:35.87" resultid="2700" heatid="6273" lane="6" entrytime="00:03:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.51" />
                    <SPLIT distance="100" swimtime="00:01:44.97" />
                    <SPLIT distance="150" swimtime="00:02:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="209" reactiontime="+108" swimtime="00:00:44.45" resultid="2701" heatid="6331" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1625" points="216" reactiontime="+100" swimtime="00:07:22.97" resultid="2702" heatid="6555" lane="1" entrytime="00:07:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.13" />
                    <SPLIT distance="100" swimtime="00:01:46.66" />
                    <SPLIT distance="150" swimtime="00:02:43.13" />
                    <SPLIT distance="200" swimtime="00:03:40.22" />
                    <SPLIT distance="250" swimtime="00:04:37.79" />
                    <SPLIT distance="300" swimtime="00:05:34.62" />
                    <SPLIT distance="350" swimtime="00:06:31.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="KU AZS Uniwersytet Wrocławski" nation="POL">
          <CONTACT city="Wrocław" email="wawrzynek77@wp.pl" name="Wawrzyńczak Karolina" phone="792777168" />
          <ATHLETES>
            <ATHLETE birthdate="1990-09-11" firstname="Karolina" gender="F" lastname="Wawrzyńczak" nation="POL" athleteid="2704">
              <RESULTS>
                <RESULT eventid="1213" points="601" reactiontime="+73" swimtime="00:00:35.30" resultid="2705" heatid="6125" lane="5" entrytime="00:00:34.80" />
                <RESULT eventid="1348" points="500" reactiontime="+86" swimtime="00:00:34.77" resultid="2706" heatid="6222" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1378" points="569" reactiontime="+70" swimtime="00:01:17.28" resultid="2707" heatid="6248" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="493" reactiontime="+87" swimtime="00:00:32.40" resultid="2708" heatid="6338" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1543" points="539" reactiontime="+71" swimtime="00:02:46.61" resultid="2709" heatid="6371" lane="4" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:21.00" />
                    <SPLIT distance="150" swimtime="00:02:04.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Astoria Bydgoszcz" nation="POL">
          <CONTACT email="sikoreczka7@o2.pl" name="Sikorska" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Krzysztof" gender="M" lastname="Kawecki" nation="POL" athleteid="2711">
              <RESULTS>
                <RESULT eventid="1092" points="681" reactiontime="+93" swimtime="00:06:24.15" resultid="2712" heatid="6489" lane="5" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:30.87" />
                    <SPLIT distance="150" swimtime="00:02:18.68" />
                    <SPLIT distance="200" swimtime="00:03:06.47" />
                    <SPLIT distance="250" swimtime="00:04:00.04" />
                    <SPLIT distance="300" swimtime="00:04:53.71" />
                    <SPLIT distance="350" swimtime="00:05:38.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="669" reactiontime="+93" swimtime="00:03:08.35" resultid="2713" heatid="6113" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                    <SPLIT distance="100" swimtime="00:01:30.04" />
                    <SPLIT distance="150" swimtime="00:02:18.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="421" reactiontime="+96" swimtime="00:03:23.05" resultid="2714" heatid="6186" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.39" />
                    <SPLIT distance="100" swimtime="00:01:35.89" />
                    <SPLIT distance="150" swimtime="00:02:27.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="521" reactiontime="+70" swimtime="00:01:23.93" resultid="2715" heatid="6255" lane="4" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="703" reactiontime="+97" swimtime="00:02:54.00" resultid="2716" heatid="6305" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:23.45" />
                    <SPLIT distance="150" swimtime="00:02:13.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="2717" heatid="6378" lane="6" entrytime="00:02:53.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BEWOP" name="Beskidzkie Wodne Ochotnicze Pogotowie Ratunkowe" nation="POL" region="KA" shortname="Beskidzkie Wodne Ochotnicze Po">
          <CONTACT city="Bielsko Biała" email="biuro@wopr.bielsko.pl" internet="http://www.wopr.bielsko.pl/" name="Eryk Gazda" phone="33-812-37-86" state="ŚLĄSK" street="1 Maja 47" zip="43-300" />
          <ATHLETES>
            <ATHLETE birthdate="1990-03-03" firstname="Magdalena" gender="F" lastname="SOLICH" nation="POL" athleteid="2720">
              <RESULTS>
                <RESULT eventid="1153" points="484" reactiontime="+82" swimtime="00:01:25.29" resultid="2721" heatid="6078" lane="4" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="492" reactiontime="+88" swimtime="00:00:41.53" resultid="2722" heatid="6199" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1595" points="468" reactiontime="+88" swimtime="00:01:30.84" resultid="2723" heatid="6509" lane="1" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-25" firstname="Roger" gender="M" lastname="ZAJĄC" nation="POL" athleteid="2724">
              <RESULTS>
                <RESULT eventid="1168" points="768" reactiontime="+64" swimtime="00:01:03.22" resultid="2725" heatid="6100" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="700" reactiontime="+68" swimtime="00:00:31.86" resultid="2726" heatid="6216" lane="6" entrytime="00:00:32.50" />
                <RESULT eventid="1528" points="784" reactiontime="+72" swimtime="00:00:24.66" resultid="2727" heatid="6354" lane="3" entrytime="00:00:28.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-03-17" firstname="Przemysław" gender="M" lastname="POBÓG-ZARZECKI" nation="POL" athleteid="2728">
              <RESULTS>
                <RESULT eventid="1333" points="432" reactiontime="+53" swimtime="00:00:39.02" resultid="2729" heatid="6205" lane="2" entrytime="00:00:45.50" />
                <RESULT eventid="1528" points="490" reactiontime="+83" swimtime="00:00:30.96" resultid="2730" heatid="6346" lane="4" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="MASTERS Białystok" nation="POL">
          <CONTACT email="epiwo@wp.pl" name="Piwowarczyk" phone="600330566" />
          <ATHLETES>
            <ATHLETE birthdate="1984-01-01" firstname="Bartosz" gender="M" lastname="Bogdanowicz" nation="POL" athleteid="2732">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="2733" heatid="6096" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="2734" heatid="6137" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1393" status="DNS" swimtime="00:00:00.00" resultid="2735" heatid="6260" lane="3" entrytime="00:01:08.00" />
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="2736" heatid="6381" lane="5" entrytime="00:02:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Joanna" gender="F" lastname="Wasilewicz" nation="POL" athleteid="2737">
              <RESULTS>
                <RESULT eventid="1257" status="DNS" swimtime="00:00:00.00" resultid="2738" heatid="6153" lane="1" entrytime="00:01:24.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="2739" heatid="6274" lane="2" entrytime="00:03:14.00" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="2740" heatid="6334" lane="1" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Mirosław" gender="M" lastname="Matusik" nation="POL" athleteid="2742">
              <RESULTS>
                <RESULT eventid="1168" points="648" reactiontime="+95" swimtime="00:01:18.60" resultid="2743" heatid="6083" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="694" reactiontime="+93" swimtime="00:03:06.01" resultid="2744" heatid="6113" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="100" swimtime="00:01:27.65" />
                    <SPLIT distance="150" swimtime="00:02:17.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="787" reactiontime="+92" swimtime="00:00:35.96" resultid="2745" heatid="6211" lane="1" entrytime="00:00:38.50" />
                <RESULT eventid="1363" points="595" swimtime="00:00:33.37" resultid="2746" heatid="6231" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1610" points="770" reactiontime="+94" swimtime="00:01:21.04" resultid="2747" heatid="6404" lane="2" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="558" reactiontime="+94" swimtime="00:05:47.57" resultid="2748" heatid="6564" lane="6" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:22.56" />
                    <SPLIT distance="150" swimtime="00:02:07.20" />
                    <SPLIT distance="200" swimtime="00:02:51.57" />
                    <SPLIT distance="250" swimtime="00:03:35.35" />
                    <SPLIT distance="300" swimtime="00:04:19.44" />
                    <SPLIT distance="350" swimtime="00:05:04.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="MOS Białystok" nation="POL">
          <CONTACT email="epiwo@wp.pl" name="Piwowarczyk" phone="600330566" />
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Marcin" gender="M" lastname="Jabłoński" nation="POL" athleteid="2750">
              <RESULTS>
                <RESULT eventid="1228" points="811" reactiontime="+57" swimtime="00:00:27.28" resultid="2751" heatid="6139" lane="2" entrytime="00:00:27.70" />
                <RESULT eventid="1272" points="863" reactiontime="+74" swimtime="00:00:51.85" resultid="2752" heatid="6180" lane="3" entrytime="00:00:52.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="782" reactiontime="+64" swimtime="00:00:59.01" resultid="2753" heatid="6262" lane="1" entrytime="00:01:01.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="804" reactiontime="+74" swimtime="00:02:12.74" resultid="2754" heatid="6311" lane="3" entrytime="00:02:12.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                    <SPLIT distance="100" swimtime="00:01:00.71" />
                    <SPLIT distance="150" swimtime="00:01:41.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="863" reactiontime="+73" swimtime="00:00:56.34" resultid="2755" heatid="6327" lane="3" entrytime="00:00:56.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="749" reactiontime="+65" swimtime="00:02:14.01" resultid="2756" heatid="6382" lane="2" entrytime="00:02:13.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:02.64" />
                    <SPLIT distance="150" swimtime="00:01:38.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="MPK Prievidza" nation="CZE">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Jozef" gender="M" lastname="Krcik" nation="CZE" athleteid="2758">
              <RESULTS>
                <RESULT eventid="1137" points="729" swimtime="00:11:07.70" resultid="2759" heatid="6452" lane="4" entrytime="00:11:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="100" swimtime="00:01:18.30" />
                    <SPLIT distance="200" swimtime="00:02:41.70" />
                    <SPLIT distance="300" swimtime="00:04:05.95" />
                    <SPLIT distance="400" swimtime="00:05:30.26" />
                    <SPLIT distance="500" swimtime="00:06:53.92" />
                    <SPLIT distance="600" swimtime="00:08:18.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="574" reactiontime="+96" swimtime="00:01:10.60" resultid="2760" heatid="6164" lane="4" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="633" reactiontime="+95" swimtime="00:02:33.49" resultid="2761" heatid="6285" lane="6" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                    <SPLIT distance="150" swimtime="00:01:54.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="696" reactiontime="+102" swimtime="00:05:22.94" resultid="2762" heatid="6565" lane="5" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:16.77" />
                    <SPLIT distance="150" swimtime="00:01:57.74" />
                    <SPLIT distance="200" swimtime="00:02:38.67" />
                    <SPLIT distance="250" swimtime="00:03:20.08" />
                    <SPLIT distance="300" swimtime="00:04:01.88" />
                    <SPLIT distance="350" swimtime="00:04:43.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Peter" gender="M" lastname="Mnasil" nation="CZE" athleteid="2763">
              <RESULTS>
                <RESULT eventid="1137" points="558" swimtime="00:12:09.90" resultid="2764" heatid="6450" lane="3" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:01:25.04" />
                    <SPLIT distance="200" swimtime="00:02:56.28" />
                    <SPLIT distance="300" swimtime="00:04:26.28" />
                    <SPLIT distance="400" swimtime="00:05:59.86" />
                    <SPLIT distance="500" swimtime="00:07:31.00" />
                    <SPLIT distance="600" swimtime="00:09:05.50" />
                    <SPLIT distance="700" swimtime="00:10:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="510" reactiontime="+105" swimtime="00:01:13.43" resultid="2765" heatid="6164" lane="3" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="609" reactiontime="+91" swimtime="00:00:39.17" resultid="2766" heatid="6207" lane="4" entrytime="00:00:43.00" />
                <RESULT eventid="1528" points="627" reactiontime="+93" swimtime="00:00:30.50" resultid="2767" heatid="6347" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1610" points="618" reactiontime="+89" swimtime="00:01:27.18" resultid="2768" heatid="6400" lane="1" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Maria" gender="F" lastname="Hausnerova" nation="CZE" athleteid="2769">
              <RESULTS>
                <RESULT eventid="1213" points="751" swimtime="00:00:42.27" resultid="2770" heatid="6122" lane="3" entrytime="00:00:42.50" />
                <RESULT eventid="1257" points="672" reactiontime="+89" swimtime="00:01:21.49" resultid="2771" heatid="6153" lane="2" entrytime="00:01:23.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="722" reactiontime="+71" swimtime="00:01:34.19" resultid="2772" heatid="6246" lane="5" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="703" reactiontime="+89" swimtime="00:00:36.15" resultid="2773" heatid="6334" lane="5" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="PVK Bratislava" nation="CZE">
          <CONTACT name="s" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Jaroslav" gender="M" lastname="Sykora" nation="CZE" athleteid="2775">
              <RESULTS>
                <RESULT eventid="1228" points="663" reactiontime="+65" swimtime="00:00:32.12" resultid="2776" heatid="6135" lane="3" entrytime="00:00:32.50" />
                <RESULT eventid="1272" points="726" reactiontime="+74" swimtime="00:00:59.42" resultid="2777" heatid="6175" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="773" reactiontime="+80" swimtime="00:00:29.04" resultid="2778" heatid="6238" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1437" points="625" reactiontime="+91" swimtime="00:02:18.41" resultid="2779" heatid="6287" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:01:05.98" />
                    <SPLIT distance="150" swimtime="00:01:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="749" reactiontime="+76" swimtime="00:00:26.89" resultid="2780" heatid="6359" lane="6" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Petr" gender="M" lastname="Soukup" nation="CZE" athleteid="2781">
              <RESULTS>
                <RESULT eventid="1272" points="748" reactiontime="+86" swimtime="00:01:00.31" resultid="2782" heatid="6174" lane="2" entrytime="00:01:00.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="656" reactiontime="+88" swimtime="00:00:35.35" resultid="2783" heatid="6214" lane="1" entrytime="00:00:34.90" />
                <RESULT eventid="1437" points="735" reactiontime="+97" swimtime="00:02:15.79" resultid="2784" heatid="6288" lane="6" entrytime="00:02:19.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:05.99" />
                    <SPLIT distance="150" swimtime="00:01:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="702" reactiontime="+84" swimtime="00:00:27.59" resultid="2785" heatid="6358" lane="4" entrytime="00:00:27.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Laura" gender="F" lastname="Majernikova" nation="CZE" athleteid="2786">
              <RESULTS>
                <RESULT eventid="1058" points="479" reactiontime="+95" swimtime="00:07:19.13" resultid="2787" heatid="6429" lane="3" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                    <SPLIT distance="100" swimtime="00:01:43.37" />
                    <SPLIT distance="150" swimtime="00:02:35.89" />
                    <SPLIT distance="200" swimtime="00:03:29.26" />
                    <SPLIT distance="250" swimtime="00:04:29.44" />
                    <SPLIT distance="300" swimtime="00:05:32.64" />
                    <SPLIT distance="350" swimtime="00:06:25.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1122" points="460" status="EXH" swimtime="00:13:18.38" resultid="2788" heatid="6443" lane="5" entrytime="00:14:19.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.46" />
                    <SPLIT distance="100" swimtime="00:01:29.45" />
                    <SPLIT distance="200" swimtime="00:03:09.27" />
                    <SPLIT distance="300" swimtime="00:04:47.81" />
                    <SPLIT distance="400" swimtime="00:06:29.90" />
                    <SPLIT distance="500" swimtime="00:08:12.91" />
                    <SPLIT distance="600" swimtime="00:09:56.31" />
                    <SPLIT distance="700" swimtime="00:11:40.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Monika" gender="F" lastname="Novakova" nation="CZE" athleteid="2789">
              <RESULTS>
                <RESULT eventid="1058" points="469" reactiontime="+90" swimtime="00:06:39.96" resultid="2790" heatid="6431" lane="6" entrytime="00:06:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:01:31.99" />
                    <SPLIT distance="150" swimtime="00:02:22.87" />
                    <SPLIT distance="200" swimtime="00:03:13.87" />
                    <SPLIT distance="250" swimtime="00:04:10.24" />
                    <SPLIT distance="300" swimtime="00:05:06.79" />
                    <SPLIT distance="350" swimtime="00:05:53.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1122" points="375" swimtime="00:12:56.88" resultid="2791" heatid="6444" lane="6" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.66" />
                    <SPLIT distance="200" swimtime="00:03:05.22" />
                    <SPLIT distance="300" swimtime="00:04:43.52" />
                    <SPLIT distance="400" swimtime="00:06:21.91" />
                    <SPLIT distance="500" swimtime="00:08:00.97" />
                    <SPLIT distance="600" swimtime="00:09:38.95" />
                    <SPLIT distance="700" swimtime="00:11:18.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="390" reactiontime="+83" swimtime="00:03:16.96" resultid="2792" heatid="6182" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.26" />
                    <SPLIT distance="100" swimtime="00:01:31.25" />
                    <SPLIT distance="150" swimtime="00:02:24.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="438" reactiontime="+91" swimtime="00:03:07.19" resultid="2793" heatid="6296" lane="1" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:29.13" />
                    <SPLIT distance="150" swimtime="00:02:24.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="357" reactiontime="+79" swimtime="00:03:15.07" resultid="2794" heatid="6368" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                    <SPLIT distance="100" swimtime="00:01:36.00" />
                    <SPLIT distance="150" swimtime="00:02:26.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+79" swimtime="00:02:05.65" resultid="2795" heatid="6496" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.40" />
                    <SPLIT distance="100" swimtime="00:01:03.28" />
                    <SPLIT distance="150" swimtime="00:01:38.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2775" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2786" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="2789" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2781" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="PHU INTER Ireneusz Nawrocki" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1989-02-25" firstname="Daniel" gender="M" lastname="Bugdol" nation="POL" athleteid="2797">
              <RESULTS>
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="4594" heatid="6456" lane="1" entrytime="00:10:00.00" />
                <RESULT eventid="1168" points="768" reactiontime="+85" swimtime="00:01:04.61" resultid="2799" heatid="6099" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="664" reactiontime="+67" swimtime="00:00:29.17" resultid="2800" heatid="6138" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1363" points="742" reactiontime="+83" swimtime="00:00:27.40" resultid="2801" heatid="6240" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="2802" heatid="6289" lane="6" entrytime="00:02:15.00" />
                <RESULT eventid="1498" points="627" reactiontime="+85" swimtime="00:01:02.68" resultid="2803" heatid="6325" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="612" reactiontime="+82" swimtime="00:00:26.28" resultid="2804" heatid="6361" lane="2" entrytime="00:00:26.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="KS Delfin Gliwice" nation="POL" region="SLA">
          <CONTACT city="Gliwice" email="ksdelfin@op.pl" name="Cupiał Jarosław" phone="605065587" state="ŚLĄSK" street="Stwosza 8/3" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Teodozja" gender="F" lastname="Gdula" nation="POL" athleteid="2806">
              <RESULTS>
                <RESULT eventid="1183" points="258" reactiontime="+132" swimtime="00:04:53.55" resultid="2807" heatid="6101" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.17" />
                    <SPLIT distance="100" swimtime="00:02:22.76" />
                    <SPLIT distance="150" swimtime="00:03:38.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="124" reactiontime="+101" swimtime="00:02:23.04" resultid="2808" heatid="6148" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="130" reactiontime="+102" swimtime="00:05:19.38" resultid="2809" heatid="6270" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.42" />
                    <SPLIT distance="100" swimtime="00:02:26.84" />
                    <SPLIT distance="150" swimtime="00:03:54.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="234" reactiontime="+105" swimtime="00:02:20.08" resultid="2810" heatid="6502" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-11-23" firstname="Jerzy" gender="M" lastname="Marciniszko" nation="POL" athleteid="2811">
              <RESULTS>
                <RESULT eventid="1198" points="182" reactiontime="+90" swimtime="00:05:25.13" resultid="2812" heatid="6108" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.17" />
                    <SPLIT distance="100" swimtime="00:02:34.24" />
                    <SPLIT distance="150" swimtime="00:04:01.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="139" reactiontime="+119" swimtime="00:01:08.01" resultid="2813" heatid="6126" lane="2" />
                <RESULT eventid="1333" points="229" reactiontime="+95" swimtime="00:00:59.08" resultid="2814" heatid="6202" lane="6" />
                <RESULT eventid="1393" points="109" reactiontime="+103" swimtime="00:02:47.36" resultid="2815" heatid="6249" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="126" reactiontime="+87" swimtime="00:00:56.28" resultid="2816" heatid="6341" lane="3" />
                <RESULT eventid="1610" points="168" reactiontime="+92" swimtime="00:02:27.36" resultid="2817" heatid="6395" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-10" firstname="Barbara" gender="F" lastname="Lipowska" nation="POL" athleteid="2818">
              <RESULTS>
                <RESULT eventid="1513" points="162" reactiontime="+104" swimtime="00:00:53.44" resultid="2819" heatid="6328" lane="5" />
                <RESULT eventid="1625" points="145" reactiontime="+104" swimtime="00:09:47.54" resultid="2820" heatid="6554" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.58" />
                    <SPLIT distance="100" swimtime="00:02:19.07" />
                    <SPLIT distance="150" swimtime="00:03:44.87" />
                    <SPLIT distance="200" swimtime="00:06:09.86" />
                    <SPLIT distance="250" swimtime="00:07:24.27" />
                    <SPLIT distance="300" swimtime="00:08:37.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Euro-Lviv" nation="UKR">
          <CONTACT city="Lviv" email="riff@mail.lviv.ua" fax="+38 032 2430304" name="Masters Swimming Club &quot;Euro-Lviv&quot;" phone="+38 067 6734796" street="Karpincya Str. 18A/3" zip="79012" />
          <ATHLETES>
            <ATHLETE birthdate="1972-09-13" firstname="Oleksandr" gender="M" lastname="Syrbu" nation="UKR" athleteid="2822">
              <RESULTS>
                <RESULT eventid="1272" points="812" reactiontime="+76" swimtime="00:00:57.25" resultid="2823" heatid="6178" lane="5" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="883" reactiontime="+77" swimtime="00:00:27.78" resultid="2824" heatid="6240" lane="4" entrytime="00:00:27.20" />
                <RESULT eventid="1528" points="800" reactiontime="+73" swimtime="00:00:26.30" resultid="2825" heatid="6364" lane="2" entrytime="00:00:25.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-05-16" firstname="Iryna" gender="F" lastname="Bura" nation="UKR" athleteid="2826">
              <RESULTS>
                <RESULT eventid="1257" points="478" reactiontime="+93" swimtime="00:01:14.24" resultid="2827" heatid="6155" lane="4" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="503" reactiontime="+94" swimtime="00:00:33.41" resultid="2828" heatid="6338" lane="1" entrytime="00:00:31.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-06-05" firstname="Mykhailo" gender="M" lastname="Shelest" nation="UKR" athleteid="2829">
              <RESULTS>
                <RESULT eventid="1228" points="548" reactiontime="+77" swimtime="00:00:38.99" resultid="2830" heatid="6132" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1333" points="662" reactiontime="+111" swimtime="00:00:38.10" resultid="2831" heatid="6211" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1610" points="668" reactiontime="+123" swimtime="00:01:24.98" resultid="2832" heatid="6403" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-08" firstname="Igor" gender="M" lastname="Rudnyk" nation="UKR" athleteid="2833">
              <RESULTS>
                <RESULT eventid="1228" points="470" reactiontime="+86" swimtime="00:00:39.37" resultid="2834" heatid="6131" lane="3" entrytime="00:00:38.50" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="2835" heatid="6346" lane="3" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-13" firstname="Bogdan" gender="M" lastname="Osidach" nation="UKR" athleteid="2836">
              <RESULTS>
                <RESULT eventid="1528" points="341" reactiontime="+93" swimtime="00:00:33.12" resultid="2837" heatid="6356" lane="6" entrytime="00:00:28.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-03" firstname="Romana" gender="F" lastname="Sirenko" nation="UKR" athleteid="2838">
              <RESULTS>
                <RESULT eventid="1153" status="DNS" swimtime="00:00:00.00" resultid="2839" heatid="6081" lane="6" entrytime="00:01:20.00" />
                <RESULT eventid="1348" status="DNS" swimtime="00:00:00.00" resultid="2840" heatid="6221" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="2841" heatid="6336" lane="3" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-07" firstname="Ruslan" gender="M" lastname="Friauf" nation="UKR" athleteid="2842">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="2843" heatid="6093" lane="1" entrytime="00:01:13.20" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="2844" heatid="6134" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="2845" heatid="6213" lane="6" entrytime="00:00:36.42" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="AZS AWF Warszawa" nation="POL">
          <CONTACT name="Gołębiowska" phone="504-794-417" />
          <ATHLETES>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="Gołębiowska" nation="POL" athleteid="2855">
              <RESULTS>
                <RESULT eventid="1153" points="924" reactiontime="+71" swimtime="00:01:06.75" resultid="2856" heatid="6082" lane="3" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. B" eventid="1348" points="960" reactiontime="+71" swimtime="00:00:29.23" resultid="2857" heatid="6223" lane="3" entrytime="00:00:29.50" />
                <RESULT comment="Rekord Polski kat. B" eventid="1422" points="858" reactiontime="+73" swimtime="00:02:11.83" resultid="2858" heatid="6277" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:04.50" />
                    <SPLIT distance="150" swimtime="00:01:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="956" reactiontime="+73" swimtime="00:01:04.93" resultid="2859" heatid="6315" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="877" reactiontime="+73" swimtime="00:00:27.76" resultid="2860" heatid="6340" lane="4" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Unlimited Triathlon Club" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1988-01-01" firstname="Marcin" gender="M" lastname="Górka" nation="POL" athleteid="2862">
              <RESULTS>
                <RESULT eventid="1228" points="641" reactiontime="+49" swimtime="00:00:29.51" resultid="2863" heatid="6139" lane="6" entrytime="00:00:29.50" />
                <RESULT eventid="1302" points="457" reactiontime="+84" swimtime="00:02:35.76" resultid="2864" heatid="6191" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                    <SPLIT distance="150" swimtime="00:01:51.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="576" reactiontime="+48" swimtime="00:01:05.35" resultid="2865" heatid="6262" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="2866" heatid="6310" lane="3" entrytime="00:02:24.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LAOLE" name="Integracyjny Miejski Klub Pływacki &quot;LAGUNA&quot; Oleśnica" nation="POL" region="DOL" shortname="Integracyjny Miejski Klub Pływ">
          <CONTACT city="Oleśnica" email="imkp.laguna@wp.pl" name="Smołuch" phone="503043978" state="DOL" street="Kopernika" zip="56-400" />
          <ATHLETES>
            <ATHLETE birthdate="1974-01-15" firstname="Artur" gender="M" lastname="Mosiak" nation="POL" athleteid="2868">
              <RESULTS>
                <RESULT eventid="1467" points="228" reactiontime="+93" swimtime="00:03:25.12" resultid="2869" heatid="6301" lane="1" entrytime="00:03:45.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:33.58" />
                    <SPLIT distance="150" swimtime="00:02:32.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-05-05" firstname="Beata" gender="F" lastname="Horbacz" nation="POL" athleteid="2870">
              <RESULTS>
                <RESULT eventid="1513" points="101" reactiontime="+125" swimtime="00:00:58.40" resultid="2871" heatid="6330" lane="4" entrytime="00:00:53.72" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-08" firstname="Adam" gender="M" lastname="Horbacz" nation="POL" athleteid="2872">
              <RESULTS>
                <RESULT eventid="1393" points="32" reactiontime="+124" swimtime="00:03:04.77" resultid="2873" heatid="6251" lane="4" entrytime="00:01:57.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Masters Kraśnik" nation="POL" region="LBL">
          <CONTACT city="Kraśnik" email="jurek@krasnik.info" internet="www.masterskrasnik.za.pl" name="Michalzyk Jerzy" phone="601698977" state="LUB" street="Żwirki i Wigury 2" zip="23-210" />
          <ATHLETES>
            <ATHLETE birthdate="1960-09-07" firstname="Andrzej" gender="M" lastname="Cis" nation="POL" athleteid="2898">
              <RESULTS>
                <RESULT eventid="1228" points="530" reactiontime="+70" swimtime="00:00:37.82" resultid="2899" heatid="6131" lane="2" entrytime="00:00:39.20" />
                <RESULT eventid="1272" points="542" reactiontime="+65" swimtime="00:01:09.77" resultid="2900" heatid="6166" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="431" swimtime="00:00:36.69" resultid="2901" heatid="6227" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1437" reactiontime="+75" status="DNS" swimtime="00:00:00.00" resultid="2902" heatid="6284" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                    <SPLIT distance="100" swimtime="00:01:16.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="553" reactiontime="+79" swimtime="00:00:30.90" resultid="2903" heatid="6350" lane="1" entrytime="00:00:31.20" />
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="2904" heatid="6375" lane="3" entrytime="00:03:19.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="2905">
              <RESULTS>
                <RESULT eventid="1168" points="320" reactiontime="+96" swimtime="00:01:39.37" resultid="2906" heatid="6083" lane="4" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="155" reactiontime="+97" swimtime="00:04:42.95" resultid="2907" heatid="6183" lane="3" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.02" />
                    <SPLIT distance="100" swimtime="00:02:14.94" />
                    <SPLIT distance="150" swimtime="00:03:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="337" reactiontime="+98" swimtime="00:00:47.71" resultid="2908" heatid="6204" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1363" points="200" swimtime="00:00:47.98" resultid="2909" heatid="6225" lane="2" entrytime="00:00:48.30" />
                <RESULT eventid="1498" points="132" reactiontime="+106" swimtime="00:02:06.15" resultid="2910" heatid="6317" lane="3" entrytime="00:01:49.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-02-09" firstname="Marcin" gender="M" lastname="Mazurek" nation="POL" athleteid="2911">
              <RESULTS>
                <RESULT eventid="1272" points="321" reactiontime="+112" swimtime="00:01:15.08" resultid="2912" heatid="6164" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="309" reactiontime="+102" swimtime="00:02:51.80" resultid="2913" heatid="6283" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:01:21.41" />
                    <SPLIT distance="150" swimtime="00:02:07.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="378" reactiontime="+99" swimtime="00:00:32.00" resultid="2914" heatid="6354" lane="1" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-27" firstname="Janusz" gender="M" lastname="Wasiuk" nation="POL" athleteid="2915">
              <RESULTS>
                <RESULT eventid="1092" points="274" reactiontime="+113" swimtime="00:08:40.13" resultid="2916" heatid="6486" lane="6" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.07" />
                    <SPLIT distance="100" swimtime="00:02:01.57" />
                    <SPLIT distance="150" swimtime="00:03:20.29" />
                    <SPLIT distance="200" swimtime="00:04:35.05" />
                    <SPLIT distance="250" swimtime="00:05:38.23" />
                    <SPLIT distance="300" swimtime="00:06:41.41" />
                    <SPLIT distance="350" swimtime="00:07:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="372" reactiontime="+118" swimtime="00:03:48.90" resultid="2917" heatid="6110" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.57" />
                    <SPLIT distance="100" swimtime="00:01:49.02" />
                    <SPLIT distance="150" swimtime="00:02:49.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="167" reactiontime="+119" swimtime="00:04:36.37" resultid="2918" heatid="6184" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.24" />
                    <SPLIT distance="100" swimtime="00:02:15.99" />
                    <SPLIT distance="150" swimtime="00:03:31.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="416" swimtime="00:00:44.46" resultid="2919" heatid="6204" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1467" points="262" reactiontime="+117" swimtime="00:04:01.76" resultid="2920" heatid="6299" lane="3" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.72" />
                    <SPLIT distance="100" swimtime="00:02:00.85" />
                    <SPLIT distance="150" swimtime="00:03:04.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="168" reactiontime="+115" swimtime="00:01:56.62" resultid="2921" heatid="6316" lane="4" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="436" reactiontime="+109" swimtime="00:01:37.96" resultid="2922" heatid="6396" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-04" firstname="Ewa" gender="F" lastname="Białosiewicz" nation="POL" athleteid="2923">
              <RESULTS>
                <RESULT eventid="1122" points="440" swimtime="00:15:01.51" resultid="2924" heatid="6443" lane="6" entrytime="00:15:00.00" />
                <RESULT eventid="1378" points="253" reactiontime="+80" swimtime="00:02:09.52" resultid="2925" heatid="6244" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="389" reactiontime="+98" swimtime="00:03:26.07" resultid="2926" heatid="6273" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                    <SPLIT distance="100" swimtime="00:01:40.97" />
                    <SPLIT distance="150" swimtime="00:02:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="366" reactiontime="+79" swimtime="00:04:19.35" resultid="2927" heatid="6368" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.51" />
                    <SPLIT distance="100" swimtime="00:02:09.36" />
                    <SPLIT distance="150" swimtime="00:03:14.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="447" reactiontime="+94" swimtime="00:07:16.13" resultid="2928" heatid="6555" lane="2" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.03" />
                    <SPLIT distance="100" swimtime="00:01:43.89" />
                    <SPLIT distance="150" swimtime="00:02:38.61" />
                    <SPLIT distance="200" swimtime="00:03:34.04" />
                    <SPLIT distance="250" swimtime="00:04:29.66" />
                    <SPLIT distance="300" swimtime="00:05:25.91" />
                    <SPLIT distance="350" swimtime="00:06:21.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" name="KS Masters Polkowice" nation="POL" region="DOL">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" state="DOL" street="Kolejowa 6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1943-11-28" firstname="Hanna" gender="F" lastname="Świder" nation="POL" athleteid="2930">
              <RESULTS>
                <RESULT eventid="1183" points="331" swimtime="00:05:12.72" resultid="2931" heatid="6102" lane="5" entrytime="00:05:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.00" />
                    <SPLIT distance="100" swimtime="00:02:28.32" />
                    <SPLIT distance="150" swimtime="00:03:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="124" swimtime="00:02:34.44" resultid="2932" heatid="6149" lane="6" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="193" swimtime="00:01:15.75" resultid="2933" heatid="6193" lane="4" entrytime="00:01:15.00" entrycourse="SCM" />
                <RESULT eventid="1422" points="138" swimtime="00:05:27.49" resultid="2934" heatid="6270" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.45" />
                    <SPLIT distance="100" swimtime="00:02:37.56" />
                    <SPLIT distance="150" swimtime="00:04:03.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="98" swimtime="00:01:15.22" resultid="2935" heatid="6329" lane="1" entrytime="00:01:12.00" entrycourse="SCM" />
                <RESULT eventid="1595" points="263" swimtime="00:02:31.68" resultid="2936" heatid="6504" lane="6" entrytime="00:02:46.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-15" firstname="Regina" gender="F" lastname="Mładszew" nation="POL" athleteid="2937">
              <RESULTS>
                <RESULT eventid="1213" points="110" reactiontime="+169" swimtime="00:01:20.18" resultid="2938" heatid="6119" lane="1" entrytime="00:01:16.00" entrycourse="SCM" />
                <RESULT eventid="1257" points="89" reactiontime="+111" swimtime="00:02:39.91" resultid="2939" heatid="6148" lane="2" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="68" reactiontime="+110" swimtime="00:01:34.46" resultid="2940" heatid="6193" lane="5" entrytime="00:01:27.00" entrycourse="SCM" />
                <RESULT eventid="1378" points="117" reactiontime="+182" swimtime="00:02:52.74" resultid="2941" heatid="6243" lane="1" entrytime="00:02:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="85" reactiontime="+108" swimtime="00:01:12.93" resultid="2942" heatid="6329" lane="5" entrytime="00:01:09.00" entrycourse="SCM" />
                <RESULT eventid="1543" points="140" reactiontime="+162" swimtime="00:06:04.00" resultid="2943" heatid="6366" lane="2" entrytime="00:06:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.47" />
                    <SPLIT distance="100" swimtime="00:02:59.70" />
                    <SPLIT distance="150" swimtime="00:04:31.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-08-16" firstname="Janina" gender="F" lastname="Zając" nation="POL" athleteid="2944">
              <RESULTS>
                <RESULT eventid="1213" points="112" reactiontime="+97" swimtime="00:01:25.13" resultid="2945" heatid="6118" lane="4" entrytime="00:01:21.00" entrycourse="SCM" />
                <RESULT eventid="1257" points="133" reactiontime="+131" swimtime="00:02:30.76" resultid="2946" heatid="6148" lane="4" entrytime="00:02:47.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="135" reactiontime="+113" swimtime="00:01:25.36" resultid="2947" heatid="6193" lane="2" entrytime="00:01:21.00" entrycourse="SCM" />
                <RESULT eventid="1378" points="142" reactiontime="+83" swimtime="00:02:57.26" resultid="2948" heatid="6242" lane="3" entrytime="00:03:08.00" entrycourse="SCM" />
                <RESULT eventid="1513" points="142" reactiontime="+111" swimtime="00:01:06.58" resultid="2949" heatid="6329" lane="2" entrytime="00:01:07.00" entrycourse="SCM" />
                <RESULT eventid="1543" points="172" reactiontime="+93" swimtime="00:06:02.49" resultid="2950" heatid="6366" lane="4" entrytime="00:06:03.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.00" />
                    <SPLIT distance="150" swimtime="00:04:34.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-05-30" firstname="Grażyna" gender="F" lastname="Grzegorzewska" nation="POL" athleteid="2951">
              <RESULTS>
                <RESULT eventid="1122" points="420" swimtime="00:16:02.50" resultid="2952" heatid="6442" lane="2" entrytime="00:15:28.00" entrycourse="SCM" />
                <RESULT eventid="1153" points="351" reactiontime="+83" swimtime="00:01:56.25" resultid="2953" heatid="6075" lane="2" entrytime="00:01:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="417" reactiontime="+84" swimtime="00:01:35.52" resultid="2954" heatid="6151" lane="6" entrytime="00:01:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="277" reactiontime="+82" swimtime="00:00:56.07" resultid="2955" heatid="6219" lane="1" entrytime="00:00:53.00" entrycourse="SCM" />
                <RESULT eventid="1422" points="390" reactiontime="+87" swimtime="00:03:41.66" resultid="2956" heatid="6273" lane="1" entrytime="00:03:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                    <SPLIT distance="100" swimtime="00:01:44.94" />
                    <SPLIT distance="150" swimtime="00:02:44.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="462" reactiontime="+86" swimtime="00:00:41.56" resultid="2957" heatid="6332" lane="1" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1625" points="414" reactiontime="+91" swimtime="00:07:41.75" resultid="2958" heatid="6555" lane="6" entrytime="00:07:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.95" />
                    <SPLIT distance="100" swimtime="00:01:48.31" />
                    <SPLIT distance="150" swimtime="00:02:48.88" />
                    <SPLIT distance="200" swimtime="00:03:48.51" />
                    <SPLIT distance="250" swimtime="00:04:48.03" />
                    <SPLIT distance="300" swimtime="00:05:47.53" />
                    <SPLIT distance="350" swimtime="00:06:47.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-10-10" firstname="Zdzisława" gender="F" lastname="Pachom" nation="POL" athleteid="2959">
              <RESULTS>
                <RESULT eventid="1153" points="66" swimtime="00:03:44.57" resultid="2960" heatid="6074" lane="2" entrytime="00:03:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="89" swimtime="00:01:38.13" resultid="2962" heatid="6193" lane="1" entrytime="00:01:33.00" entrycourse="SCM" />
                <RESULT eventid="1348" points="52" swimtime="00:01:45.00" resultid="2963" heatid="6218" lane="1" entrytime="00:01:41.00" entrycourse="SCM" />
                <RESULT eventid="1513" points="95" swimtime="00:01:16.01" resultid="2964" heatid="6328" lane="2" entrytime="00:01:37.00" entrycourse="SCM" />
                <RESULT eventid="1595" points="102" swimtime="00:03:27.68" resultid="2965" heatid="6503" lane="4" entrytime="00:03:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:42.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="111" swimtime="00:07:28.93" resultid="6539" heatid="6101" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:44.47" />
                    <SPLIT distance="100" swimtime="00:03:37.15" />
                    <SPLIT distance="150" swimtime="00:05:31.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-10-02" firstname="Emilia" gender="F" lastname="Kawula" nation="POL" athleteid="2966">
              <RESULTS>
                <RESULT eventid="1257" points="92" swimtime="00:03:10.70" resultid="2968" heatid="6148" lane="3" entrytime="00:02:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="103" swimtime="00:01:34.82" resultid="2969" heatid="6193" lane="6" entrytime="00:01:34.00" entrycourse="SCM" />
                <RESULT eventid="1513" points="97" swimtime="00:01:21.83" resultid="2970" heatid="6329" lane="6" entrytime="00:01:12.00" entrycourse="SCM" />
                <RESULT eventid="1595" points="99" swimtime="00:03:35.11" resultid="2971" heatid="6503" lane="2" entrytime="00:03:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:43.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="131" swimtime="00:07:25.62" resultid="6547" heatid="6107" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.49" />
                    <SPLIT distance="100" swimtime="00:03:36.86" />
                    <SPLIT distance="150" swimtime="00:05:31.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-02" firstname="Wiesław" gender="M" lastname="Zając" nation="POL" athleteid="2972">
              <RESULTS>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="2973" heatid="6108" lane="4" entrytime="00:04:53.00" entrycourse="SCM" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="2974" heatid="6160" lane="6" entrytime="00:01:54.00" entrycourse="SCM" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="2975" heatid="6202" lane="4" entrytime="00:01:04.00" entrycourse="SCM" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="2976" heatid="6278" lane="4" entrytime="00:04:27.00" entrycourse="SCM" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="2977" heatid="6342" lane="4" entrytime="00:00:48.00" entrycourse="SCM" />
                <RESULT eventid="1610" status="DNS" swimtime="00:00:00.00" resultid="2978" heatid="6395" lane="4" entrytime="00:02:18.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-05-26" firstname="Zygmunt" gender="M" lastname="Pawlaczek" nation="POL" athleteid="2979">
              <RESULTS>
                <RESULT eventid="1137" points="272" swimtime="00:15:36.62" resultid="2980" heatid="6447" lane="2" entrytime="00:17:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                    <SPLIT distance="100" swimtime="00:01:36.50" />
                    <SPLIT distance="200" swimtime="00:03:29.11" />
                    <SPLIT distance="300" swimtime="00:05:28.01" />
                    <SPLIT distance="400" swimtime="00:07:30.02" />
                    <SPLIT distance="500" swimtime="00:09:32.08" />
                    <SPLIT distance="600" swimtime="00:11:36.08" />
                    <SPLIT distance="700" swimtime="00:13:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z2" eventid="1168" reactiontime="+110" status="DSQ" swimtime="00:01:35.67" resultid="2981" heatid="6086" lane="5" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="463" reactiontime="+98" swimtime="00:01:20.60" resultid="2982" heatid="6162" lane="6" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="387" reactiontime="+119" swimtime="00:03:13.70" resultid="2983" heatid="6279" lane="3" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                    <SPLIT distance="100" swimtime="00:01:28.17" />
                    <SPLIT distance="150" swimtime="00:02:20.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="319" reactiontime="+103" swimtime="00:07:11.80" resultid="2984" heatid="6561" lane="2" entrytime="00:06:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:01:30.25" />
                    <SPLIT distance="150" swimtime="00:02:24.55" />
                    <SPLIT distance="200" swimtime="00:03:20.62" />
                    <SPLIT distance="250" swimtime="00:04:17.04" />
                    <SPLIT distance="300" swimtime="00:05:14.64" />
                    <SPLIT distance="350" swimtime="00:06:13.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-04-23" firstname="Bogdan" gender="M" lastname="Jawor" nation="POL" athleteid="2985">
              <RESULTS>
                <RESULT eventid="1137" points="282" swimtime="00:17:15.88" resultid="2986" heatid="6447" lane="3" entrytime="00:16:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.03" />
                    <SPLIT distance="100" swimtime="00:01:47.85" />
                    <SPLIT distance="200" swimtime="00:03:53.39" />
                    <SPLIT distance="300" swimtime="00:05:57.17" />
                    <SPLIT distance="400" swimtime="00:08:03.35" />
                    <SPLIT distance="500" swimtime="00:10:06.59" />
                    <SPLIT distance="600" swimtime="00:12:10.06" />
                    <SPLIT distance="700" swimtime="00:14:12.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="268" reactiontime="+98" swimtime="00:01:57.12" resultid="2987" heatid="6083" lane="3" entrytime="00:01:53.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="311" reactiontime="+93" swimtime="00:04:32.19" resultid="2988" heatid="6109" lane="6" entrytime="00:04:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.04" />
                    <SPLIT distance="100" swimtime="00:02:12.28" />
                    <SPLIT distance="150" swimtime="00:03:25.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="318" reactiontime="+81" swimtime="00:00:52.98" resultid="2989" heatid="6203" lane="4" entrytime="00:00:54.00" entrycourse="SCM" />
                <RESULT eventid="1437" points="291" reactiontime="+101" swimtime="00:03:44.18" resultid="2990" heatid="6279" lane="6" entrytime="00:03:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.84" />
                    <SPLIT distance="100" swimtime="00:01:47.14" />
                    <SPLIT distance="150" swimtime="00:02:47.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="239" reactiontime="+86" swimtime="00:04:40.99" resultid="2991" heatid="6372" lane="4" entrytime="00:04:44.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.89" />
                    <SPLIT distance="100" swimtime="00:02:18.23" />
                    <SPLIT distance="150" swimtime="00:03:29.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="288" reactiontime="+103" swimtime="00:02:03.28" resultid="2992" heatid="6396" lane="1" entrytime="00:01:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-03" firstname="Ewa" gender="F" lastname="Puchalska" nation="POL" athleteid="2993">
              <RESULTS>
                <RESULT eventid="1183" points="192" reactiontime="+98" swimtime="00:05:09.13" resultid="2994" heatid="6102" lane="2" entrytime="00:05:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.46" />
                    <SPLIT distance="100" swimtime="00:02:31.14" />
                    <SPLIT distance="150" swimtime="00:03:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="123" reactiontime="+167" swimtime="00:01:09.50" resultid="2995" heatid="6119" lane="5" entrytime="00:01:07.00" entrycourse="SCM" />
                <RESULT eventid="1318" points="232" reactiontime="+86" swimtime="00:01:01.64" resultid="2996" heatid="6193" lane="3" entrytime="00:01:05.00" entrycourse="SCM" />
                <RESULT eventid="1378" points="114" reactiontime="+104" swimtime="00:02:39.10" resultid="2997" heatid="6243" lane="5" entrytime="00:02:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="103" reactiontime="+97" swimtime="00:01:02.12" resultid="2998" heatid="6330" lane="5" entrytime="00:00:57.00" entrycourse="SCM" />
                <RESULT eventid="1595" points="214" reactiontime="+89" swimtime="00:02:19.22" resultid="2999" heatid="6504" lane="1" entrytime="00:02:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-06-21" firstname="Bogdan" gender="M" lastname="Puchalski" nation="POL" athleteid="3000">
              <RESULTS>
                <RESULT eventid="1168" points="400" reactiontime="+85" swimtime="00:01:32.29" resultid="3001" heatid="6087" lane="5" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="341" reactiontime="+70" swimtime="00:00:45.65" resultid="3002" heatid="6130" lane="5" entrytime="00:00:43.00" entrycourse="SCM" />
                <RESULT eventid="1333" points="423" reactiontime="+83" swimtime="00:00:44.21" resultid="3003" heatid="6207" lane="5" entrytime="00:00:44.00" entrycourse="SCM" />
                <RESULT eventid="1363" points="342" reactiontime="+90" swimtime="00:00:40.14" resultid="3004" heatid="6227" lane="6" entrytime="00:00:39.00" entrycourse="SCM" />
                <RESULT eventid="1528" points="478" reactiontime="+84" swimtime="00:00:33.38" resultid="3005" heatid="6347" lane="2" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1610" points="460" reactiontime="+93" swimtime="00:01:36.20" resultid="3006" heatid="6398" lane="3" entrytime="00:01:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-02" firstname="Zenon" gender="M" lastname="Wilk" nation="POL" athleteid="3007">
              <RESULTS>
                <RESULT eventid="1168" points="73" reactiontime="+115" swimtime="00:02:51.93" resultid="3008" heatid="6083" lane="5" entrytime="00:02:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="122" reactiontime="+69" swimtime="00:01:07.38" resultid="3009" heatid="6127" lane="6" entrytime="00:01:02.00" entrycourse="SCM" />
                <RESULT eventid="1363" points="40" reactiontime="+120" swimtime="00:01:28.54" resultid="3010" heatid="6224" lane="5" entrytime="00:01:15.00" entrycourse="SCM" />
                <RESULT eventid="1393" points="107" reactiontime="+77" swimtime="00:02:34.80" resultid="3011" heatid="6250" lane="4" entrytime="00:02:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="133" reactiontime="+68" swimtime="00:05:16.96" resultid="3012" heatid="6372" lane="2" entrytime="00:05:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.66" />
                    <SPLIT distance="100" swimtime="00:02:33.20" />
                    <SPLIT distance="150" swimtime="00:03:56.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-02" firstname="Pavlo" gender="M" lastname="Vechirko" nation="POL" athleteid="3013">
              <RESULTS>
                <RESULT eventid="1198" points="591" reactiontime="+106" swimtime="00:02:59.13" resultid="3014" heatid="6114" lane="6" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:25.03" />
                    <SPLIT distance="150" swimtime="00:02:10.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="520" reactiontime="+72" swimtime="00:01:15.49" resultid="3015" heatid="6258" lane="4" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="578" reactiontime="+78" swimtime="00:02:42.65" resultid="3016" heatid="6380" lane="6" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="150" swimtime="00:01:59.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="536" reactiontime="+166" swimtime="00:01:22.70" resultid="3017" heatid="6402" lane="4" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+78" swimtime="00:02:42.38" resultid="3020" heatid="6521" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                    <SPLIT distance="100" swimtime="00:01:27.97" />
                    <SPLIT distance="150" swimtime="00:02:07.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3013" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="2985" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3000" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="2979" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="O4 - przedwczesny start." eventid="1415" status="DSQ" swimtime="00:02:28.12" resultid="3021" heatid="6529" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:01:52.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2985" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="3013" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="3000" number="3" reactiontime="+45" status="DSQ" />
                    <RELAYPOSITION athleteid="2979" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1243" reactiontime="+167" swimtime="00:04:23.48" resultid="3018" heatid="6519" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.83" />
                    <SPLIT distance="100" swimtime="00:02:20.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2937" number="1" reactiontime="+167" />
                    <RELAYPOSITION athleteid="2993" number="2" reactiontime="+15" />
                    <RELAYPOSITION athleteid="2951" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2944" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1408" reactiontime="+110" swimtime="00:04:07.93" resultid="3019" heatid="6527" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.28" />
                    <SPLIT distance="100" swimtime="00:02:23.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2937" number="1" reactiontime="+110" />
                    <RELAYPOSITION athleteid="2944" number="2" reactiontime="-109" />
                    <RELAYPOSITION athleteid="2993" number="3" reactiontime="+92" />
                    <RELAYPOSITION athleteid="2951" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+180" swimtime="00:04:11.09" resultid="3023" heatid="6535" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2937" number="1" reactiontime="+180" />
                    <RELAYPOSITION athleteid="2944" number="2" />
                    <RELAYPOSITION athleteid="2985" number="3" />
                    <RELAYPOSITION athleteid="2979" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+73" swimtime="00:03:04.67" resultid="3022" heatid="6535" lane="4">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:22.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3013" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="2993" number="2" />
                    <RELAYPOSITION athleteid="3000" number="3" />
                    <RELAYPOSITION athleteid="2951" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="K.S. niezrzeszeni.pl" nation="POL">
          <CONTACT email="niezrzeszenipl@mail.com" internet="niezezwszeni.pl" name="Wawer Matylda Katarzyna" phone="501701359" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="3038">
              <RESULTS>
                <RESULT eventid="1092" points="325" reactiontime="+109" swimtime="00:07:39.79" resultid="3039" heatid="6486" lane="2" entrytime="00:08:25.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.97" />
                    <SPLIT distance="100" swimtime="00:01:48.01" />
                    <SPLIT distance="150" swimtime="00:03:44.40" />
                    <SPLIT distance="200" swimtime="00:04:48.33" />
                    <SPLIT distance="250" swimtime="00:05:56.57" />
                    <SPLIT distance="300" swimtime="00:06:51.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="377" reactiontime="+121" swimtime="00:01:30.67" resultid="3040" heatid="6086" lane="4" entrytime="00:01:31.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="417" reactiontime="+63" swimtime="00:00:40.98" resultid="3041" heatid="6130" lane="3" entrytime="00:00:40.26" />
                <RESULT eventid="1393" points="402" reactiontime="+63" swimtime="00:01:31.03" resultid="3042" heatid="6254" lane="2" entrytime="00:01:29.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="436" reactiontime="+57" swimtime="00:03:16.38" resultid="3043" heatid="6376" lane="6" entrytime="00:03:17.54">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:27.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-08-26" firstname="Małgorzata" gender="F" lastname="Piechura" nation="POL" athleteid="3044">
              <RESULTS>
                <RESULT eventid="1122" points="142" swimtime="00:17:53.56" resultid="3045" heatid="6441" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.46" />
                    <SPLIT distance="100" swimtime="00:01:57.42" />
                    <SPLIT distance="200" swimtime="00:04:09.64" />
                    <SPLIT distance="300" swimtime="00:06:27.83" />
                    <SPLIT distance="400" swimtime="00:08:46.54" />
                    <SPLIT distance="500" swimtime="00:11:04.13" />
                    <SPLIT distance="600" swimtime="00:13:21.62" />
                    <SPLIT distance="700" swimtime="00:15:40.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="269" reactiontime="+119" swimtime="00:04:08.25" resultid="3046" heatid="6103" lane="3" entrytime="00:04:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.91" />
                    <SPLIT distance="100" swimtime="00:02:00.74" />
                    <SPLIT distance="150" swimtime="00:03:06.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="154" reactiontime="+111" swimtime="00:01:47.65" resultid="3047" heatid="6149" lane="4" entrytime="00:01:54.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="252" reactiontime="+114" swimtime="00:00:52.95" resultid="3048" heatid="6195" lane="4" entrytime="00:00:52.80" />
                <RESULT eventid="1422" points="137" reactiontime="+119" swimtime="00:04:03.58" resultid="3049" heatid="6271" lane="5" entrytime="00:04:15.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.12" />
                    <SPLIT distance="100" swimtime="00:01:55.42" />
                    <SPLIT distance="150" swimtime="00:02:59.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="162" reactiontime="+112" swimtime="00:00:49.09" resultid="3050" heatid="6330" lane="3" entrytime="00:00:48.89" />
                <RESULT eventid="1625" points="143" reactiontime="+116" swimtime="00:08:31.00" resultid="3051" heatid="6554" lane="2" entrytime="00:08:45.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.53" />
                    <SPLIT distance="100" swimtime="00:01:56.94" />
                    <SPLIT distance="150" swimtime="00:03:01.46" />
                    <SPLIT distance="200" swimtime="00:04:05.64" />
                    <SPLIT distance="250" swimtime="00:05:11.68" />
                    <SPLIT distance="300" swimtime="00:06:19.07" />
                    <SPLIT distance="350" swimtime="00:07:28.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-14" firstname="Andrzej" gender="M" lastname="Miński" nation="POL" athleteid="3052">
              <RESULTS>
                <RESULT eventid="1137" points="409" swimtime="00:13:29.68" resultid="3053" heatid="6450" lane="6" entrytime="00:12:38.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:01:30.84" />
                    <SPLIT distance="200" swimtime="00:03:09.34" />
                    <SPLIT distance="300" swimtime="00:04:50.72" />
                    <SPLIT distance="400" swimtime="00:06:33.10" />
                    <SPLIT distance="500" swimtime="00:08:16.57" />
                    <SPLIT distance="600" swimtime="00:10:01.32" />
                    <SPLIT distance="700" swimtime="00:11:47.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="437" reactiontime="+107" swimtime="00:03:37.06" resultid="3054" heatid="6111" lane="3" entrytime="00:03:29.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.48" />
                    <SPLIT distance="100" swimtime="00:01:44.26" />
                    <SPLIT distance="150" swimtime="00:02:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="370" reactiontime="+110" swimtime="00:01:21.74" resultid="3055" heatid="6161" lane="4" entrytime="00:01:20.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="414" swimtime="00:00:44.53" resultid="3056" heatid="6207" lane="2" entrytime="00:00:43.84" />
                <RESULT eventid="1437" points="383" reactiontime="+107" swimtime="00:03:01.45" resultid="3057" heatid="6281" lane="1" entrytime="00:02:59.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:26.36" />
                    <SPLIT distance="150" swimtime="00:02:14.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="425" reactiontime="+105" swimtime="00:01:38.81" resultid="3058" heatid="6398" lane="5" entrytime="00:01:38.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="409" reactiontime="+104" swimtime="00:06:25.67" resultid="3059" heatid="6562" lane="3" entrytime="00:06:17.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="100" swimtime="00:01:30.84" />
                    <SPLIT distance="150" swimtime="00:02:20.10" />
                    <SPLIT distance="200" swimtime="00:03:09.13" />
                    <SPLIT distance="250" swimtime="00:03:58.42" />
                    <SPLIT distance="300" swimtime="00:04:48.30" />
                    <SPLIT distance="350" swimtime="00:05:38.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="SGGW Warszawa" nation="POL">
          <CONTACT city="Warszawa" email="olszewski_krzysiek@o2.pl" name="Olszewski" street="Nowoursynowska 166" />
          <ATHLETES>
            <ATHLETE birthdate="1989-07-28" firstname="Krzysztof" gender="M" lastname="Olszewski" nation="POL" athleteid="3061">
              <RESULTS>
                <RESULT comment="G5" eventid="1168" reactiontime="+75" status="DSQ" swimtime="00:01:08.08" resultid="3062" heatid="6098" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="561" reactiontime="+76" swimtime="00:00:59.84" resultid="3063" heatid="6176" lane="5" entrytime="00:00:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="617" reactiontime="+74" swimtime="00:00:33.27" resultid="3064" heatid="6215" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="1467" points="561" reactiontime="+77" swimtime="00:02:29.67" resultid="3065" heatid="6308" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:10.13" />
                    <SPLIT distance="150" swimtime="00:01:52.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="614" reactiontime="+77" swimtime="00:00:26.26" resultid="3066" heatid="6363" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1610" points="594" reactiontime="+75" swimtime="00:01:13.93" resultid="3067" heatid="6407" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Legia Warszawa" nation="POL">
          <CONTACT email="janek@plywanielegia.pl" internet="www.plywanielegia.pl" name="Drzewiński" phone="600826305" />
          <ATHLETES>
            <ATHLETE birthdate="1986-08-28" firstname="Krzesimir" gender="M" lastname="Sieczych" nation="POL" athleteid="3069">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="3070" heatid="6094" lane="2" entrytime="00:01:12.00" />
                <RESULT eventid="1363" status="DNS" swimtime="00:00:00.00" resultid="3071" heatid="6235" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3072" heatid="6359" lane="4" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-16" firstname="Maciej" gender="M" lastname="Drzewiński" nation="POL" athleteid="3093">
              <RESULTS>
                <RESULT eventid="1363" status="DNS" swimtime="00:00:00.00" resultid="3094" heatid="6238" lane="1" entrytime="00:00:29.20" />
                <RESULT eventid="1528" points="697" reactiontime="+70" swimtime="00:00:26.02" resultid="3095" heatid="6362" lane="5" entrytime="00:00:26.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-09" firstname="Tomasz" gender="M" lastname="Drzewiński" nation="POL" athleteid="3096">
              <RESULTS>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3097" heatid="6205" lane="5" entrytime="00:00:45.80" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3098" heatid="6349" lane="3" entrytime="00:00:31.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-03-09" firstname="Łukasz" gender="M" lastname="Drzewiński" nation="POL" athleteid="3099">
              <RESULTS>
                <RESULT eventid="1168" points="875" reactiontime="+73" swimtime="00:01:00.54" resultid="3100" heatid="6100" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="884" reactiontime="+75" swimtime="00:00:26.42" resultid="3101" heatid="6241" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1498" points="886" reactiontime="+78" swimtime="00:00:57.82" resultid="3102" heatid="6327" lane="4" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-26" firstname="Tomasz" gender="M" lastname="Wilczęga" nation="POL" athleteid="3103">
              <RESULTS>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3104" heatid="6362" lane="4" entrytime="00:00:26.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-24" firstname="Marcin" gender="M" lastname="Wilczęga" nation="POL" athleteid="3105">
              <RESULTS>
                <RESULT eventid="1528" points="628" reactiontime="+74" swimtime="00:00:26.93" resultid="3106" heatid="6362" lane="2" entrytime="00:00:26.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-27" firstname="Jan" gender="M" lastname="Peńsko" nation="POL" athleteid="3107">
              <RESULTS>
                <RESULT eventid="1168" points="833" reactiontime="+82" swimtime="00:01:01.53" resultid="3108" heatid="6100" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="806" reactiontime="+67" swimtime="00:00:28.09" resultid="3109" heatid="6139" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="1393" points="766" reactiontime="+72" swimtime="00:01:01.42" resultid="3110" heatid="6262" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="862" reactiontime="+85" swimtime="00:00:58.35" resultid="3112" heatid="6327" lane="2" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="819" reactiontime="+77" swimtime="00:02:13.52" resultid="3113" heatid="6382" lane="5" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:06.48" />
                    <SPLIT distance="150" swimtime="00:01:40.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-12" firstname="Krzysztof" gender="M" lastname="Spyra" nation="POL" athleteid="3114">
              <RESULTS>
                <RESULT eventid="1437" points="565" reactiontime="+97" swimtime="00:02:20.50" resultid="3115" heatid="6284" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:08.17" />
                    <SPLIT distance="150" swimtime="00:01:44.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="530" reactiontime="+85" swimtime="00:00:28.60" resultid="3116" heatid="6354" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1640" points="522" reactiontime="+91" swimtime="00:05:04.81" resultid="3117" heatid="6566" lane="2" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:09.83" />
                    <SPLIT distance="150" swimtime="00:01:48.28" />
                    <SPLIT distance="200" swimtime="00:02:27.01" />
                    <SPLIT distance="250" swimtime="00:03:06.93" />
                    <SPLIT distance="300" swimtime="00:03:46.64" />
                    <SPLIT distance="350" swimtime="00:04:26.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-06-08" firstname="Maciej" gender="M" lastname="Grzelak" nation="POL" athleteid="3118">
              <RESULTS>
                <RESULT eventid="1092" points="360" reactiontime="+86" swimtime="00:06:52.35" resultid="3119" heatid="6488" lane="1" entrytime="00:06:56.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                    <SPLIT distance="100" swimtime="00:01:24.00" />
                    <SPLIT distance="150" swimtime="00:02:24.89" />
                    <SPLIT distance="200" swimtime="00:03:25.21" />
                    <SPLIT distance="250" swimtime="00:04:22.13" />
                    <SPLIT distance="300" swimtime="00:05:21.07" />
                    <SPLIT distance="350" swimtime="00:06:07.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="464" reactiontime="+77" swimtime="00:01:19.70" resultid="3120" heatid="6089" lane="3" entrytime="00:01:20.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="301" reactiontime="+74" swimtime="00:03:14.60" resultid="3121" heatid="6186" lane="5" entrytime="00:03:20.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:01:25.20" />
                    <SPLIT distance="150" swimtime="00:02:20.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="496" reactiontime="+79" swimtime="00:00:33.68" resultid="3122" heatid="6228" lane="4" entrytime="00:00:35.61" />
                <RESULT eventid="1467" points="445" reactiontime="+81" swimtime="00:02:58.63" resultid="3123" heatid="6303" lane="3" entrytime="00:03:09.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:27.29" />
                    <SPLIT distance="150" swimtime="00:02:18.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="425" reactiontime="+79" swimtime="00:01:17.98" resultid="3124" heatid="6321" lane="1" entrytime="00:01:19.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="424" reactiontime="+81" swimtime="00:01:29.42" resultid="3125" heatid="6398" lane="1" entrytime="00:01:38.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+67" swimtime="00:01:58.68" resultid="3073" heatid="6526" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                    <SPLIT distance="150" swimtime="00:01:32.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3107" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3096" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3099" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3093" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1415" reactiontime="+73" swimtime="00:01:41.50" resultid="3074" heatid="6534" lane="3" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                    <SPLIT distance="100" swimtime="00:00:52.17" />
                    <SPLIT distance="150" swimtime="00:01:16.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3105" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3093" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="3099" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3107" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+77" swimtime="00:02:11.76" resultid="3075" heatid="6526" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="150" swimtime="00:01:43.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3103" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3105" number="2" reactiontime="+17" />
                    <RELAYPOSITION athleteid="3118" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3114" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1415" reactiontime="+76" swimtime="00:02:07.17" resultid="3076" heatid="6534" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                    <SPLIT distance="100" swimtime="00:00:59.10" />
                    <SPLIT distance="150" swimtime="00:01:38.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3103" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3118" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3096" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="3114" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Delfin Gdynia" nation="POL">
          <CONTACT name="s" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Jakub" gender="M" lastname="Mańczak" nation="POL" athleteid="3127">
              <RESULTS>
                <RESULT eventid="1302" points="523" reactiontime="+82" swimtime="00:02:41.84" resultid="3128" heatid="6190" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:15.55" />
                    <SPLIT distance="150" swimtime="00:02:00.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="772" reactiontime="+76" swimtime="00:00:29.06" resultid="3129" heatid="6237" lane="4" entrytime="00:00:29.70" />
                <RESULT eventid="1498" points="628" reactiontime="+78" swimtime="00:01:08.48" resultid="3130" heatid="6324" lane="3" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="704" reactiontime="+77" swimtime="00:00:27.45" resultid="3131" heatid="6358" lane="2" entrytime="00:00:27.60" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MACHE" name="Masters Chełm" nation="POL">
          <CONTACT city="Chełm" email="elzbietadz@gmail.com" name="Dziwisz  Elżbieta" phone="660429651" state="LUBEL" street="Lubelska 139 D/13" zip="22-100" />
          <ATHLETES>
            <ATHLETE birthdate="1954-01-01" firstname="Elżbieta" gender="F" lastname="Dziwisz" nation="POL" athleteid="3133">
              <RESULTS>
                <RESULT eventid="1183" points="258" reactiontime="+98" swimtime="00:04:58.08" resultid="3134" heatid="6103" lane="5" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.86" />
                    <SPLIT distance="100" swimtime="00:02:24.63" />
                    <SPLIT distance="150" swimtime="00:03:41.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="254" reactiontime="+89" swimtime="00:00:58.47" resultid="3135" heatid="6119" lane="4" entrytime="00:01:02.00" />
                <RESULT eventid="1318" points="253" reactiontime="+100" swimtime="00:01:00.77" resultid="3136" heatid="6194" lane="6" entrytime="00:00:58.00" />
                <RESULT eventid="1378" points="260" reactiontime="+83" swimtime="00:02:08.45" resultid="3137" heatid="6244" lane="5" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="185" reactiontime="+98" swimtime="00:00:54.35" resultid="3138" heatid="6330" lane="2" entrytime="00:00:54.00" />
                <RESULT eventid="1595" points="255" reactiontime="+98" swimtime="00:02:17.64" resultid="3139" heatid="6505" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Hanna" gender="F" lastname="Wepa" nation="POL" athleteid="3140">
              <RESULTS>
                <RESULT eventid="1122" points="102" swimtime="00:22:26.69" resultid="3141" heatid="6441" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.29" />
                    <SPLIT distance="100" swimtime="00:02:36.23" />
                    <SPLIT distance="150" swimtime="00:03:58.41" />
                    <SPLIT distance="200" swimtime="00:05:20.61" />
                    <SPLIT distance="250" swimtime="00:06:42.34" />
                    <SPLIT distance="300" swimtime="00:08:07.06" />
                    <SPLIT distance="350" swimtime="00:09:32.55" />
                    <SPLIT distance="400" swimtime="00:10:55.42" />
                    <SPLIT distance="450" swimtime="00:12:21.64" />
                    <SPLIT distance="500" swimtime="00:13:48.16" />
                    <SPLIT distance="550" swimtime="00:15:16.10" />
                    <SPLIT distance="600" swimtime="00:16:42.53" />
                    <SPLIT distance="650" swimtime="00:18:10.64" />
                    <SPLIT distance="700" swimtime="00:19:37.32" />
                    <SPLIT distance="750" swimtime="00:21:01.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="203" reactiontime="+119" swimtime="00:05:03.60" resultid="3142" heatid="6103" lane="6" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.49" />
                    <SPLIT distance="100" swimtime="00:02:27.40" />
                    <SPLIT distance="150" swimtime="00:03:46.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="88" reactiontime="+121" swimtime="00:02:26.22" resultid="3143" heatid="6149" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="194" reactiontime="+134" swimtime="00:01:05.41" resultid="3144" heatid="6194" lane="4" entrytime="00:00:55.00" />
                <RESULT eventid="1422" points="99" reactiontime="+135" swimtime="00:05:09.21" resultid="3145" heatid="6271" lane="1" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.28" />
                    <SPLIT distance="100" swimtime="00:02:27.87" />
                    <SPLIT distance="150" swimtime="00:03:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="171" reactiontime="+116" swimtime="00:02:30.17" resultid="3146" heatid="6504" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="89" reactiontime="+125" swimtime="00:11:30.04" resultid="3147" heatid="6554" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.53" />
                    <SPLIT distance="100" swimtime="00:02:41.20" />
                    <SPLIT distance="150" swimtime="00:04:06.10" />
                    <SPLIT distance="200" swimtime="00:05:35.84" />
                    <SPLIT distance="250" swimtime="00:07:07.79" />
                    <SPLIT distance="300" swimtime="00:08:36.36" />
                    <SPLIT distance="350" swimtime="00:10:03.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Wiesław" gender="M" lastname="Wepa" nation="POL" athleteid="3148">
              <RESULTS>
                <RESULT eventid="1137" points="221" swimtime="00:16:33.86" resultid="3149" heatid="6446" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.05" />
                    <SPLIT distance="100" swimtime="00:01:43.59" />
                    <SPLIT distance="200" swimtime="00:03:38.66" />
                    <SPLIT distance="300" swimtime="00:05:39.59" />
                    <SPLIT distance="400" swimtime="00:07:48.58" />
                    <SPLIT distance="500" swimtime="00:10:02.34" />
                    <SPLIT distance="600" swimtime="00:12:10.94" />
                    <SPLIT distance="700" swimtime="00:14:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="251" reactiontime="+98" swimtime="00:01:47.76" resultid="3150" heatid="6084" lane="3" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="336" reactiontime="+98" swimtime="00:03:56.93" resultid="3151" heatid="6109" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.58" />
                    <SPLIT distance="100" swimtime="00:01:55.55" />
                    <SPLIT distance="150" swimtime="00:02:56.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="340" reactiontime="+95" swimtime="00:00:47.58" resultid="3152" heatid="6202" lane="5" entrytime="00:01:44.00" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="3153" heatid="6301" lane="6" entrytime="00:03:50.00" />
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="3154" heatid="6373" lane="4" entrytime="00:04:00.00" />
                <RESULT eventid="1610" points="327" reactiontime="+101" swimtime="00:01:47.81" resultid="3155" heatid="6397" lane="5" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Janusz" gender="M" lastname="Golik" nation="POL" athleteid="3156">
              <RESULTS>
                <RESULT eventid="1198" points="543" reactiontime="+109" swimtime="00:03:58.85" resultid="3157" heatid="6110" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.19" />
                    <SPLIT distance="100" swimtime="00:01:58.25" />
                    <SPLIT distance="150" swimtime="00:03:00.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="386" reactiontime="+113" swimtime="00:04:25.84" resultid="3158" heatid="6184" lane="3" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.76" />
                    <SPLIT distance="100" swimtime="00:02:11.81" />
                    <SPLIT distance="150" swimtime="00:03:19.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="622" reactiontime="+112" swimtime="00:00:44.77" resultid="3159" heatid="6208" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1363" points="383" reactiontime="+100" swimtime="00:00:46.94" resultid="3160" heatid="6225" lane="4" entrytime="00:00:47.00" />
                <RESULT eventid="1498" points="355" reactiontime="+102" swimtime="00:01:53.70" resultid="3161" heatid="6317" lane="5" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="535" reactiontime="+113" swimtime="00:01:47.82" resultid="3162" heatid="6397" lane="1" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1107" swimtime="00:03:29.22" resultid="3163" heatid="6494" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.24" />
                    <SPLIT distance="100" swimtime="00:01:58.42" />
                    <SPLIT distance="150" swimtime="00:02:40.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3133" number="1" />
                    <RELAYPOSITION athleteid="3140" number="2" />
                    <RELAYPOSITION athleteid="3156" number="3" />
                    <RELAYPOSITION athleteid="3148" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1588" reactiontime="+80" swimtime="00:03:48.53" resultid="3164" heatid="6535" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.18" />
                    <SPLIT distance="100" swimtime="00:02:14.33" />
                    <SPLIT distance="150" swimtime="00:03:04.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3133" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3140" number="2" reactiontime="-105" />
                    <RELAYPOSITION athleteid="3156" number="3" />
                    <RELAYPOSITION athleteid="3148" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MASGOR" name="MASTERS Gorzów Wlkp." nation="POL" region="LBS">
          <CONTACT city="Gorzów Wlkp." email="woycek@poczta.onet.pl" name="Wojciechowicz Marek" phone="602891603" state="LUB" street="Ogińskiego 97/7" zip="66-400" />
          <ATHLETES>
            <ATHLETE birthdate="1970-12-12" firstname="Marek" gender="M" lastname="Wojciechowicz" nation="POL" license="MWOJ" athleteid="3166">
              <RESULTS>
                <RESULT eventid="1137" points="523" swimtime="00:10:42.24" resultid="3167" heatid="6453" lane="1" entrytime="00:11:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:10.44" />
                    <SPLIT distance="200" swimtime="00:02:28.89" />
                    <SPLIT distance="300" swimtime="00:03:50.51" />
                    <SPLIT distance="400" swimtime="00:05:12.51" />
                    <SPLIT distance="500" swimtime="00:06:35.01" />
                    <SPLIT distance="600" swimtime="00:07:58.51" />
                    <SPLIT distance="700" swimtime="00:09:22.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="700" reactiontime="+87" swimtime="00:01:00.15" resultid="3168" heatid="6173" lane="2" entrytime="00:01:01.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="647" reactiontime="+76" swimtime="00:02:16.81" resultid="3169" heatid="6285" lane="3" entrytime="00:02:30.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                    <SPLIT distance="100" swimtime="00:01:03.92" />
                    <SPLIT distance="150" swimtime="00:01:40.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="695" reactiontime="+78" swimtime="00:00:27.56" resultid="3170" heatid="6358" lane="3" entrytime="00:00:27.57" entrycourse="SCM" />
                <RESULT eventid="1640" points="566" reactiontime="+92" swimtime="00:05:03.61" resultid="3171" heatid="6566" lane="4" entrytime="00:05:18.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:09.28" />
                    <SPLIT distance="150" swimtime="00:01:48.01" />
                    <SPLIT distance="200" swimtime="00:02:27.41" />
                    <SPLIT distance="250" swimtime="00:03:06.98" />
                    <SPLIT distance="300" swimtime="00:03:46.82" />
                    <SPLIT distance="350" swimtime="00:04:26.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-20" firstname="Artur" gender="M" lastname="Rutkowski" nation="POL" license="ARUT" athleteid="3178">
              <RESULTS>
                <RESULT eventid="1092" points="490" reactiontime="+87" swimtime="00:06:01.80" resultid="3179" heatid="6488" lane="4" entrytime="00:06:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:01:18.51" />
                    <SPLIT distance="150" swimtime="00:02:06.42" />
                    <SPLIT distance="200" swimtime="00:02:53.39" />
                    <SPLIT distance="250" swimtime="00:03:46.16" />
                    <SPLIT distance="300" swimtime="00:04:39.95" />
                    <SPLIT distance="350" swimtime="00:05:22.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="433" reactiontime="+87" swimtime="00:02:51.63" resultid="3180" heatid="6188" lane="3" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:17.02" />
                    <SPLIT distance="150" swimtime="00:02:04.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="457" reactiontime="+86" swimtime="00:02:42.77" resultid="3181" heatid="6306" lane="1" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:16.23" />
                    <SPLIT distance="150" swimtime="00:02:04.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="467" reactiontime="+90" swimtime="00:01:13.53" resultid="3182" heatid="6322" lane="2" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" license="MLAS" athleteid="3183">
              <RESULTS>
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="3184" heatid="6448" lane="2" entrytime="00:14:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Orka Mastes Radlin" nation="POL">
          <CONTACT email="otelom.080966interia.pl" name="otlik marian" phone="530556313" />
          <ATHLETES>
            <ATHLETE birthdate="1940-08-10" firstname="JAN" gender="M" lastname="KLAPSIA" nation="POL" athleteid="3196">
              <RESULTS>
                <RESULT eventid="1228" points="135" swimtime="00:01:14.33" resultid="3197" heatid="6126" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="1272" points="58" reactiontime="+124" swimtime="00:02:52.52" resultid="3198" heatid="6159" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="153" swimtime="00:01:11.44" resultid="3199" heatid="6202" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="1528" points="93" reactiontime="+125" swimtime="00:01:06.53" resultid="3201" heatid="6342" lane="1" entrytime="00:01:10.00" />
                <RESULT eventid="1610" points="115" reactiontime="+114" swimtime="00:02:59.98" resultid="3202" heatid="6395" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="102" reactiontime="+98" swimtime="00:03:00.62" resultid="6546" heatid="6249" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-16" firstname="BUGLA" gender="M" lastname="RUDOLF" nation="POL" athleteid="3203">
              <RESULTS>
                <RESULT eventid="1092" points="417" reactiontime="+109" swimtime="00:08:49.78" resultid="3204" heatid="6485" lane="3" entrytime="00:08:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.06" />
                    <SPLIT distance="100" swimtime="00:02:02.47" />
                    <SPLIT distance="150" swimtime="00:03:10.20" />
                    <SPLIT distance="200" swimtime="00:04:19.77" />
                    <SPLIT distance="250" swimtime="00:05:29.08" />
                    <SPLIT distance="300" swimtime="00:06:39.01" />
                    <SPLIT distance="350" swimtime="00:07:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="323" reactiontime="+81" swimtime="00:00:55.67" resultid="3205" heatid="6128" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1302" points="419" reactiontime="+106" swimtime="00:04:18.61" resultid="3206" heatid="6185" lane="1" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.35" />
                    <SPLIT distance="100" swimtime="00:02:05.61" />
                    <SPLIT distance="150" swimtime="00:03:11.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="294" reactiontime="+99" swimtime="00:00:51.29" resultid="3207" heatid="6225" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1467" points="438" reactiontime="+108" swimtime="00:04:04.58" resultid="3208" heatid="6300" lane="5" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.25" />
                    <SPLIT distance="100" swimtime="00:01:57.79" />
                    <SPLIT distance="150" swimtime="00:03:03.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="326" reactiontime="+94" swimtime="00:01:56.96" resultid="3209" heatid="6317" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="389" reactiontime="+94" swimtime="00:04:13.71" resultid="3210" heatid="6373" lane="1" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.26" />
                    <SPLIT distance="100" swimtime="00:02:03.20" />
                    <SPLIT distance="150" swimtime="00:03:08.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-07" firstname="LEON" gender="M" lastname="IRCZYK" nation="POL" athleteid="3211">
              <RESULTS>
                <RESULT eventid="1092" points="352" reactiontime="+126" swimtime="00:08:13.12" resultid="3212" heatid="6486" lane="5" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.56" />
                    <SPLIT distance="100" swimtime="00:02:04.30" />
                    <SPLIT distance="150" swimtime="00:03:07.69" />
                    <SPLIT distance="200" swimtime="00:05:15.82" />
                    <SPLIT distance="250" swimtime="00:06:17.26" />
                    <SPLIT distance="300" swimtime="00:07:16.34" />
                    <SPLIT distance="350" swimtime="00:08:19.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="453" reactiontime="+138" swimtime="00:03:49.76" resultid="3213" heatid="6109" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.19" />
                    <SPLIT distance="100" swimtime="00:01:52.96" />
                    <SPLIT distance="150" swimtime="00:02:51.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="213" reactiontime="+113" swimtime="00:04:31.27" resultid="3214" heatid="6184" lane="4" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.55" />
                    <SPLIT distance="100" swimtime="00:02:12.61" />
                    <SPLIT distance="150" swimtime="00:03:22.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="258" reactiontime="+122" swimtime="00:03:41.60" resultid="3215" heatid="6279" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                    <SPLIT distance="100" swimtime="00:01:42.00" />
                    <SPLIT distance="150" swimtime="00:02:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="323" reactiontime="+145" swimtime="00:03:54.60" resultid="3216" heatid="6300" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.25" />
                    <SPLIT distance="100" swimtime="00:02:59.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="151" reactiontime="+111" swimtime="00:02:11.36" resultid="3217" heatid="6317" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="238" reactiontime="+121" swimtime="00:07:56.10" resultid="3218" heatid="6561" lane="6" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.19" />
                    <SPLIT distance="100" swimtime="00:01:52.04" />
                    <SPLIT distance="150" swimtime="00:02:52.94" />
                    <SPLIT distance="200" swimtime="00:03:54.20" />
                    <SPLIT distance="250" swimtime="00:04:56.13" />
                    <SPLIT distance="300" swimtime="00:05:57.32" />
                    <SPLIT distance="350" swimtime="00:06:57.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="JERZY" gender="M" lastname="CIECIOR" nation="POL" athleteid="3219">
              <RESULTS>
                <RESULT eventid="1137" points="485" swimtime="00:12:44.85" resultid="3220" heatid="6451" lane="6" entrytime="00:12:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.95" />
                    <SPLIT distance="200" swimtime="00:03:01.59" />
                    <SPLIT distance="300" swimtime="00:04:38.92" />
                    <SPLIT distance="400" swimtime="00:06:16.12" />
                    <SPLIT distance="500" swimtime="00:07:54.26" />
                    <SPLIT distance="600" swimtime="00:09:31.35" />
                    <SPLIT distance="700" swimtime="00:11:11.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="448" reactiontime="+88" swimtime="00:01:28.83" resultid="3221" heatid="6088" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="509" reactiontime="+53" swimtime="00:00:39.95" resultid="3222" heatid="6131" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1393" points="432" reactiontime="+61" swimtime="00:01:29.38" resultid="3223" heatid="6254" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="3224" heatid="6282" lane="5" entrytime="00:02:45.00" />
                <RESULT eventid="1498" points="426" reactiontime="+74" swimtime="00:01:25.50" resultid="3225" heatid="6320" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="429" reactiontime="+80" swimtime="00:03:19.57" resultid="3226" heatid="6375" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:35.63" />
                    <SPLIT distance="150" swimtime="00:02:28.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-08-08" firstname="SŁAWOMIR" gender="M" lastname="SZUREK" nation="POL" athleteid="3227">
              <RESULTS>
                <RESULT eventid="1092" points="366" reactiontime="+92" swimtime="00:06:50.14" resultid="3228" heatid="6487" lane="4" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:01:28.27" />
                    <SPLIT distance="150" swimtime="00:03:17.61" />
                    <SPLIT distance="200" swimtime="00:04:14.14" />
                    <SPLIT distance="250" swimtime="00:05:13.19" />
                    <SPLIT distance="300" swimtime="00:06:02.15" />
                    <SPLIT distance="350" swimtime="00:06:50.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="406" reactiontime="+90" swimtime="00:01:23.33" resultid="3229" heatid="6091" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="389" reactiontime="+89" swimtime="00:01:13.13" resultid="3230" heatid="6167" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="426" reactiontime="+91" swimtime="00:00:35.43" resultid="3231" heatid="6229" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1467" points="398" reactiontime="+84" swimtime="00:03:05.30" resultid="3232" heatid="6303" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:29.51" />
                    <SPLIT distance="150" swimtime="00:02:22.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="443" reactiontime="+95" swimtime="00:00:32.02" resultid="3233" heatid="6351" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1640" points="372" reactiontime="+90" swimtime="00:05:49.24" resultid="3234" heatid="6564" lane="1" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:20.01" />
                    <SPLIT distance="150" swimtime="00:02:04.17" />
                    <SPLIT distance="200" swimtime="00:02:49.13" />
                    <SPLIT distance="250" swimtime="00:03:34.43" />
                    <SPLIT distance="300" swimtime="00:04:20.34" />
                    <SPLIT distance="350" swimtime="00:05:06.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-24" firstname="PIOTR" gender="M" lastname="SOBIK" nation="POL" athleteid="3235">
              <RESULTS>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3236" heatid="6205" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1363" points="343" reactiontime="+93" swimtime="00:00:36.06" resultid="3237" heatid="6228" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1498" points="263" reactiontime="+105" swimtime="00:01:26.92" resultid="3238" heatid="6318" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="227" reactiontime="+107" swimtime="00:00:37.79" resultid="3239" heatid="6343" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1610" status="DNS" swimtime="00:00:00.00" resultid="3240" heatid="6401" lane="1" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-09" firstname="TOMASZ" gender="M" lastname="ŻURCZAK" nation="POL" athleteid="3241">
              <RESULTS>
                <RESULT eventid="1137" points="317" swimtime="00:12:38.80" resultid="3242" heatid="6449" lane="3" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:25.58" />
                    <SPLIT distance="200" swimtime="00:03:00.24" />
                    <SPLIT distance="300" swimtime="00:04:34.81" />
                    <SPLIT distance="400" swimtime="00:06:11.66" />
                    <SPLIT distance="500" swimtime="00:07:48.16" />
                    <SPLIT distance="600" swimtime="00:09:25.44" />
                    <SPLIT distance="700" swimtime="00:11:01.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="389" reactiontime="+94" swimtime="00:03:25.87" resultid="3243" heatid="6108" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                    <SPLIT distance="100" swimtime="00:01:36.02" />
                    <SPLIT distance="150" swimtime="00:02:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="3244" heatid="6161" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3245" heatid="6210" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="3246" heatid="6281" lane="6" entrytime="00:03:00.00" />
                <RESULT eventid="1528" points="361" reactiontime="+93" swimtime="00:00:34.29" resultid="3247" heatid="6345" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1610" points="383" reactiontime="+90" swimtime="00:01:32.48" resultid="3248" heatid="6399" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-09" firstname="MARIAN" gender="M" lastname="OTLIK" nation="POL" athleteid="3249">
              <RESULTS>
                <RESULT eventid="1092" points="382" reactiontime="+100" swimtime="00:06:58.44" resultid="3250" heatid="6487" lane="3" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:32.83" />
                    <SPLIT distance="200" swimtime="00:03:25.01" />
                    <SPLIT distance="300" swimtime="00:05:24.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="465" reactiontime="+76" swimtime="00:01:22.05" resultid="3251" heatid="6089" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="486" reactiontime="+77" swimtime="00:01:09.64" resultid="3252" heatid="6165" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="432" swimtime="00:00:36.22" resultid="3253" heatid="6228" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1467" points="401" reactiontime="+85" swimtime="00:03:09.48" resultid="3254" heatid="6303" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                    <SPLIT distance="100" swimtime="00:01:30.22" />
                    <SPLIT distance="150" swimtime="00:02:26.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="523" reactiontime="+72" swimtime="00:00:30.43" resultid="3255" heatid="6348" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1610" points="373" reactiontime="+68" swimtime="00:01:35.50" resultid="3256" heatid="6399" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-06-25" firstname="EWA" gender="F" lastname="ADAMCZYK" nation="POL" athleteid="3257">
              <RESULTS>
                <RESULT eventid="1183" points="329" reactiontime="+104" swimtime="00:03:56.51" resultid="3258" heatid="6104" lane="3" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.77" />
                    <SPLIT distance="100" swimtime="00:01:50.99" />
                    <SPLIT distance="150" swimtime="00:02:55.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="381" reactiontime="+91" swimtime="00:00:46.91" resultid="3260" heatid="6198" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1422" points="223" reactiontime="+98" swimtime="00:03:34.20" resultid="3261" heatid="6272" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.29" />
                    <SPLIT distance="100" swimtime="00:01:43.97" />
                    <SPLIT distance="150" swimtime="00:02:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="342" reactiontime="+84" swimtime="00:00:38.86" resultid="3262" heatid="6332" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1595" points="387" reactiontime="+98" swimtime="00:01:43.10" resultid="3263" heatid="6507" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="248" reactiontime="+87" swimtime="00:01:33.75" resultid="6549" heatid="6151" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-08-06" firstname="RENATA" gender="F" lastname="MACIOŃCZYK" nation="POL" athleteid="3264">
              <RESULTS>
                <RESULT eventid="1183" points="305" reactiontime="+88" swimtime="00:03:58.27" resultid="3265" heatid="6104" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.69" />
                    <SPLIT distance="100" swimtime="00:01:54.49" />
                    <SPLIT distance="150" swimtime="00:02:57.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="277" reactiontime="+90" swimtime="00:01:28.44" resultid="3266" heatid="6152" lane="4" entrytime="00:01:25.00" />
                <RESULT eventid="1318" points="341" reactiontime="+65" swimtime="00:00:47.87" resultid="3267" heatid="6196" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="3268" heatid="6271" lane="4" entrytime="00:04:00.00" />
                <RESULT eventid="1513" points="350" reactiontime="+90" swimtime="00:00:38.00" resultid="3269" heatid="6335" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1595" points="344" reactiontime="+82" swimtime="00:01:45.80" resultid="3270" heatid="6506" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+78" swimtime="00:03:25.82" resultid="6025" heatid="6521" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="100" swimtime="00:01:52.57" />
                    <SPLIT distance="150" swimtime="00:02:48.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3196" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3203" number="2" reactiontime="+96" />
                    <RELAYPOSITION athleteid="3211" number="3" reactiontime="-161" />
                    <RELAYPOSITION athleteid="3219" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+78" swimtime="00:02:29.93" resultid="6026" heatid="6521" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:23.84" />
                    <SPLIT distance="150" swimtime="00:02:00.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3227" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3241" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="3235" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3249" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+88" swimtime="00:02:12.07" resultid="6027" heatid="6529" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:06.87" />
                    <SPLIT distance="150" swimtime="00:01:40.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3235" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="3249" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="3241" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3227" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+105" status="DNS" swimtime="00:00:00.00" resultid="3271" heatid="6529" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3196" number="1" reactiontime="+105" />
                    <RELAYPOSITION athleteid="3211" number="2" reactiontime="+94" />
                    <RELAYPOSITION athleteid="3219" number="3" />
                    <RELAYPOSITION athleteid="3203" number="4" reactiontime="+79" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+59" swimtime="00:02:40.34" resultid="3272" heatid="6535" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:01:27.25" />
                    <SPLIT distance="150" swimtime="00:02:02.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3219" number="1" reactiontime="+59" />
                    <RELAYPOSITION athleteid="3257" number="2" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3227" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="3264" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="MOSiR Piekary Śląskie" nation="POL">
          <CONTACT name="Szymik" />
          <ATHLETES>
            <ATHLETE birthdate="1986-03-07" firstname="Bartosz" gender="M" lastname="Szymik" nation="POL" athleteid="3276">
              <RESULTS>
                <RESULT eventid="1198" points="519" reactiontime="+98" swimtime="00:02:56.65" resultid="3277" heatid="6115" lane="1" entrytime="00:02:57.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                    <SPLIT distance="100" swimtime="00:01:24.37" />
                    <SPLIT distance="150" swimtime="00:02:10.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="378" reactiontime="+74" swimtime="00:02:52.76" resultid="3278" heatid="6378" lane="1" entrytime="00:02:50.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                    <SPLIT distance="100" swimtime="00:01:23.03" />
                    <SPLIT distance="150" swimtime="00:02:08.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="523" reactiontime="+91" swimtime="00:01:18.43" resultid="3279" heatid="6404" lane="3" entrytime="00:01:20.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01103" name="MTP Lublinianka" nation="POL" region="LU">
          <CONTACT name="Mazurek" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-26" firstname="Jarosław" gender="M" lastname="Mazurek" nation="POL" license="S01103200003" athleteid="3281">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. B" eventid="1137" points="738" swimtime="00:09:11.68" resultid="3282" heatid="6446" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                    <SPLIT distance="100" swimtime="00:01:00.54" />
                    <SPLIT distance="200" swimtime="00:02:06.55" />
                    <SPLIT distance="300" swimtime="00:03:13.87" />
                    <SPLIT distance="400" swimtime="00:04:23.48" />
                    <SPLIT distance="500" swimtime="00:05:35.31" />
                    <SPLIT distance="600" swimtime="00:06:48.52" />
                    <SPLIT distance="700" swimtime="00:08:01.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="888" reactiontime="+68" swimtime="00:00:27.16" resultid="3283" heatid="6139" lane="3" entrytime="00:00:26.25" />
                <RESULT eventid="1272" points="817" reactiontime="+79" swimtime="00:00:54.18" resultid="3284" heatid="6180" lane="4" entrytime="00:00:53.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="898" reactiontime="+69" swimtime="00:00:58.73" resultid="3285" heatid="6262" lane="3" entrytime="00:00:57.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="840" reactiontime="+76" swimtime="00:01:58.32" resultid="3286" heatid="6292" lane="3" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.61" />
                    <SPLIT distance="100" swimtime="00:00:57.84" />
                    <SPLIT distance="150" swimtime="00:01:28.35" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. B" eventid="1558" points="911" reactiontime="+71" swimtime="00:02:10.39" resultid="3287" heatid="6382" lane="3" entrytime="00:02:06.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                    <SPLIT distance="100" swimtime="00:01:01.68" />
                    <SPLIT distance="150" swimtime="00:01:35.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="TMT &quot;Water Knights&quot; Zabierzów" nation="POL">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1976-01-01" firstname="Artur" gender="M" lastname="Czerwiec" nation="POL" athleteid="3302">
              <RESULTS>
                <RESULT eventid="1137" points="583" swimtime="00:10:16.51" resultid="3303" heatid="6455" lane="3" entrytime="00:10:10.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:07.05" />
                    <SPLIT distance="200" swimtime="00:02:20.74" />
                    <SPLIT distance="300" swimtime="00:03:37.38" />
                    <SPLIT distance="400" swimtime="00:04:56.51" />
                    <SPLIT distance="500" swimtime="00:06:16.54" />
                    <SPLIT distance="600" swimtime="00:07:38.03" />
                    <SPLIT distance="700" swimtime="00:08:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="648" reactiontime="+80" swimtime="00:00:59.42" resultid="3304" heatid="6177" lane="5" entrytime="00:00:58.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="678" reactiontime="+84" swimtime="00:02:12.24" resultid="3305" heatid="6291" lane="4" entrytime="00:02:08.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:03.69" />
                    <SPLIT distance="150" swimtime="00:01:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="633" reactiontime="+81" swimtime="00:00:26.95" resultid="3306" heatid="6360" lane="3" entrytime="00:00:26.79" />
                <RESULT eventid="1640" points="617" reactiontime="+86" swimtime="00:04:48.25" resultid="3307" heatid="6569" lane="6" entrytime="00:04:45.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="100" swimtime="00:01:07.82" />
                    <SPLIT distance="150" swimtime="00:01:44.60" />
                    <SPLIT distance="200" swimtime="00:02:21.79" />
                    <SPLIT distance="250" swimtime="00:02:58.54" />
                    <SPLIT distance="300" swimtime="00:03:35.36" />
                    <SPLIT distance="350" swimtime="00:04:12.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Grzegorz" gender="M" lastname="Mytnik" nation="POL" athleteid="3864">
              <RESULTS>
                <RESULT eventid="1137" points="367" swimtime="00:12:02.68" resultid="3865" heatid="6451" lane="1" entrytime="00:12:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:13.24" />
                    <SPLIT distance="200" swimtime="00:02:44.35" />
                    <SPLIT distance="300" swimtime="00:04:15.35" />
                    <SPLIT distance="400" swimtime="00:05:48.20" />
                    <SPLIT distance="500" swimtime="00:07:21.37" />
                    <SPLIT distance="600" swimtime="00:08:56.32" />
                    <SPLIT distance="700" swimtime="00:10:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="406" reactiontime="+101" swimtime="00:05:39.05" resultid="3866" heatid="6566" lane="5" entrytime="00:05:20.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:16.78" />
                    <SPLIT distance="150" swimtime="00:01:57.78" />
                    <SPLIT distance="200" swimtime="00:02:41.87" />
                    <SPLIT distance="350" swimtime="00:04:55.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Pływalnia Oceanik Ostrzeszów" nation="POL">
          <CONTACT city="Ostrzeszów" name="Burghardt Nina" phone="660945504" street="Kąpielowa 4a" zip="63-500" />
          <ATHLETES>
            <ATHLETE birthdate="1986-06-21" firstname="Nina" gender="F" lastname="Burghardt" nation="POL" athleteid="3309">
              <RESULTS>
                <RESULT eventid="1153" points="669" reactiontime="+77" swimtime="00:01:14.96" resultid="3310" heatid="6081" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. A" eventid="1213" points="835" reactiontime="+64" swimtime="00:00:32.33" resultid="3311" heatid="6125" lane="3" entrytime="00:00:32.60" />
                <RESULT eventid="1318" points="806" reactiontime="+76" swimtime="00:00:36.62" resultid="3312" heatid="6201" lane="1" entrytime="00:00:37.50" />
                <RESULT eventid="1348" points="744" reactiontime="+75" swimtime="00:00:32.16" resultid="3313" heatid="6223" lane="1" entrytime="00:00:32.30" />
                <RESULT eventid="1378" status="DNS" swimtime="00:00:00.00" resultid="3314" heatid="6248" lane="3" entrytime="00:01:13.50" />
                <RESULT eventid="1513" points="651" reactiontime="+75" swimtime="00:00:30.45" resultid="3315" heatid="6340" lane="6" entrytime="00:00:29.90" />
                <RESULT eventid="1595" points="674" reactiontime="+74" swimtime="00:01:20.64" resultid="3316" heatid="6510" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Wodnik Radom" nation="POL">
          <CONTACT name="Pajdzik" />
          <ATHLETES>
            <ATHLETE birthdate="1960-01-06" firstname="Andrzej" gender="M" lastname="Średnicki" nation="POL" athleteid="3318">
              <RESULTS>
                <RESULT eventid="1137" points="503" swimtime="00:11:52.82" resultid="3319" heatid="6453" lane="3" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                    <SPLIT distance="100" swimtime="00:01:21.32" />
                    <SPLIT distance="200" swimtime="00:02:49.13" />
                    <SPLIT distance="300" swimtime="00:04:19.46" />
                    <SPLIT distance="400" swimtime="00:05:50.22" />
                    <SPLIT distance="500" swimtime="00:07:22.32" />
                    <SPLIT distance="600" swimtime="00:08:53.86" />
                    <SPLIT distance="700" swimtime="00:10:25.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="3320" heatid="6114" lane="4" entrytime="00:03:00.00" />
                <RESULT eventid="1272" points="557" reactiontime="+76" swimtime="00:01:09.12" resultid="3321" heatid="6170" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="3322" heatid="6286" lane="1" entrytime="00:02:30.00" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="3323" heatid="6306" lane="5" entrytime="00:02:50.00" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3324" heatid="6354" lane="5" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PIKON" name="UKS &quot;Piątka&quot; Konstantynów Łódzki" nation="POL" region="LOD" shortname="UKS &quot;Piątka&quot; Konstantynów Łódz">
          <CONTACT email="tomaszkotus@tlen.pl" name="Kotus Tomasz" phone="603820602" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Marcin" gender="M" lastname="Grabarczyk" nation="POL" athleteid="3327">
              <RESULTS>
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="3328" heatid="6455" lane="2" entrytime="00:10:17.77" />
                <RESULT eventid="1168" points="568" reactiontime="+79" swimtime="00:01:10.36" resultid="3329" heatid="6091" lane="3" entrytime="00:01:17.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="457" reactiontime="+81" swimtime="00:03:02.41" resultid="3330" heatid="6116" lane="4" entrytime="00:02:47.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                    <SPLIT distance="100" swimtime="00:01:23.53" />
                    <SPLIT distance="150" swimtime="00:02:11.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="424" reactiontime="+68" swimtime="00:01:15.39" resultid="3331" heatid="6255" lane="3" entrytime="00:01:21.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="561" reactiontime="+82" swimtime="00:02:35.96" resultid="3332" heatid="6308" lane="3" entrytime="00:02:37.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:59.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="3333" heatid="6378" lane="3" entrytime="00:02:47.77" />
                <RESULT eventid="1640" points="538" reactiontime="+80" swimtime="00:04:55.71" resultid="3334" heatid="6567" lane="2" entrytime="00:04:57.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:07.93" />
                    <SPLIT distance="150" swimtime="00:01:43.66" />
                    <SPLIT distance="200" swimtime="00:02:20.65" />
                    <SPLIT distance="250" swimtime="00:02:58.26" />
                    <SPLIT distance="300" swimtime="00:03:37.58" />
                    <SPLIT distance="350" swimtime="00:04:16.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-02" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="3335">
              <RESULTS>
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="3336" heatid="6452" lane="5" entrytime="00:11:45.00" />
                <RESULT eventid="1198" points="412" reactiontime="+97" swimtime="00:03:08.85" resultid="3337" heatid="6116" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:28.35" />
                    <SPLIT distance="150" swimtime="00:02:19.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="416" reactiontime="+73" swimtime="00:00:34.96" resultid="3338" heatid="6138" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1333" points="467" swimtime="00:00:37.95" resultid="3339" heatid="6216" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1393" points="391" reactiontime="+79" swimtime="00:01:17.45" resultid="3340" heatid="6259" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="385" reactiontime="+64" swimtime="00:02:53.73" resultid="3341" heatid="6379" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:02:08.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="484" reactiontime="+96" swimtime="00:01:22.60" resultid="3342" heatid="6402" lane="6" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-02" firstname="Jakub" gender="M" lastname="Gryczyński" nation="POL" athleteid="3343">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="3344" heatid="6090" lane="4" entrytime="00:01:20.00" />
                <RESULT eventid="1333" points="453" reactiontime="+89" swimtime="00:00:38.35" resultid="3345" heatid="6211" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1610" points="416" reactiontime="+80" swimtime="00:01:26.89" resultid="3346" heatid="6401" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-05" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" athleteid="3347">
              <RESULTS>
                <RESULT eventid="1272" points="539" reactiontime="+97" swimtime="00:01:02.21" resultid="3348" heatid="6172" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="529" reactiontime="+96" swimtime="00:00:31.22" resultid="3349" heatid="6231" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1528" points="646" reactiontime="+89" swimtime="00:00:26.68" resultid="3350" heatid="6357" lane="2" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-05" firstname="Witold" gender="M" lastname="Pietrowski" nation="POL" athleteid="3351">
              <RESULTS>
                <RESULT eventid="1272" points="414" reactiontime="+80" swimtime="00:01:07.95" resultid="3352" heatid="6167" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="531" reactiontime="+87" swimtime="00:00:31.19" resultid="3353" heatid="6231" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3354" heatid="6352" lane="2" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-09" firstname="Damian" gender="M" lastname="Karkusiński" nation="POL" athleteid="3355">
              <RESULTS>
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="3356" heatid="6134" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="3357" heatid="6167" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="1393" status="DNS" swimtime="00:00:00.00" resultid="3358" heatid="6259" lane="6" entrytime="00:01:14.00" />
                <RESULT comment="O4 - przedwczesny start." eventid="1528" reactiontime="+51" status="DSQ" swimtime="00:00:31.16" resultid="3359" heatid="6352" lane="4" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-03" firstname="Rafał" gender="M" lastname="Trudnos" nation="POL" athleteid="3360">
              <RESULTS>
                <RESULT eventid="1168" points="473" reactiontime="+79" swimtime="00:01:14.77" resultid="3361" heatid="6095" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="651" reactiontime="+81" swimtime="00:00:33.99" resultid="3362" heatid="6216" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1363" points="567" reactiontime="+79" swimtime="00:00:30.51" resultid="3363" heatid="6236" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1610" points="585" reactiontime="+79" swimtime="00:01:17.57" resultid="3364" heatid="6407" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-09-09" firstname="Igor" gender="M" lastname="Olejarczyk" nation="POL" athleteid="3365">
              <RESULTS>
                <RESULT eventid="1272" points="568" reactiontime="+83" swimtime="00:01:01.13" resultid="3366" heatid="6175" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="620" reactiontime="+88" swimtime="00:00:29.62" resultid="3367" heatid="6236" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1437" points="366" reactiontime="+93" swimtime="00:02:36.04" resultid="3368" heatid="6286" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:13.03" />
                    <SPLIT distance="150" swimtime="00:01:54.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="514" reactiontime="+83" swimtime="00:01:09.53" resultid="3369" heatid="6324" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="660" reactiontime="+79" swimtime="00:00:26.49" resultid="3370" heatid="6357" lane="5" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-03" firstname="Łukasz" gender="M" lastname="Raj" nation="POL" athleteid="3371">
              <RESULTS>
                <RESULT eventid="1092" points="337" reactiontime="+105" swimtime="00:06:34.70" resultid="3372" heatid="6490" lane="1" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:26.02" />
                    <SPLIT distance="150" swimtime="00:02:20.10" />
                    <SPLIT distance="200" swimtime="00:03:12.20" />
                    <SPLIT distance="250" swimtime="00:04:07.66" />
                    <SPLIT distance="300" swimtime="00:05:02.64" />
                    <SPLIT distance="350" swimtime="00:05:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="3373" heatid="6171" lane="4" entrytime="00:01:03.00" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3374" heatid="6213" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1528" points="413" reactiontime="+82" swimtime="00:00:30.96" resultid="3375" heatid="6354" lane="6" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-08" firstname="Kornel" gender="M" lastname="Pintara" nation="POL" athleteid="3376">
              <RESULTS>
                <RESULT eventid="1272" points="544" reactiontime="+91" swimtime="00:01:02.04" resultid="3377" heatid="6170" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="526" swimtime="00:00:31.28" resultid="3378" heatid="6234" lane="2" entrytime="00:00:30.86" />
                <RESULT eventid="1437" points="434" reactiontime="+91" swimtime="00:02:27.40" resultid="3379" heatid="6286" lane="2" entrytime="00:02:25.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:13.17" />
                    <SPLIT distance="150" swimtime="00:01:51.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="554" reactiontime="+83" swimtime="00:00:28.08" resultid="3380" heatid="6358" lane="6" entrytime="00:00:27.86" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" athleteid="3381">
              <RESULTS>
                <RESULT eventid="1137" points="529" swimtime="00:10:36.68" resultid="3382" heatid="6456" lane="5" entrytime="00:09:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:09.53" />
                    <SPLIT distance="200" swimtime="00:02:25.47" />
                    <SPLIT distance="300" swimtime="00:03:44.54" />
                    <SPLIT distance="400" swimtime="00:05:05.15" />
                    <SPLIT distance="500" swimtime="00:06:27.17" />
                    <SPLIT distance="600" swimtime="00:07:50.94" />
                    <SPLIT distance="700" swimtime="00:09:15.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="523" reactiontime="+85" swimtime="00:01:12.46" resultid="3383" heatid="6099" lane="4" entrytime="00:01:03.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="598" reactiontime="+79" swimtime="00:01:01.02" resultid="3384" heatid="6176" lane="1" entrytime="00:00:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="613" reactiontime="+79" swimtime="00:00:29.59" resultid="3385" heatid="6237" lane="6" entrytime="00:00:29.99" />
                <RESULT eventid="1437" points="604" reactiontime="+80" swimtime="00:02:17.44" resultid="3386" heatid="6291" lane="5" entrytime="00:02:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:05.49" />
                    <SPLIT distance="150" swimtime="00:01:41.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="595" reactiontime="+78" swimtime="00:00:27.52" resultid="3387" heatid="6357" lane="4" entrytime="00:00:27.99" />
                <RESULT eventid="1640" points="596" reactiontime="+79" swimtime="00:04:51.57" resultid="3388" heatid="6568" lane="3" entrytime="00:04:49.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="100" swimtime="00:01:09.61" />
                    <SPLIT distance="150" swimtime="00:01:46.17" />
                    <SPLIT distance="200" swimtime="00:02:23.84" />
                    <SPLIT distance="250" swimtime="00:03:01.24" />
                    <SPLIT distance="300" swimtime="00:03:38.94" />
                    <SPLIT distance="350" swimtime="00:04:16.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-04" firstname="Jakub" gender="M" lastname="Sidorowicz" nation="POL" athleteid="3389">
              <RESULTS>
                <RESULT eventid="1198" points="284" reactiontime="+82" swimtime="00:03:35.91" resultid="3390" heatid="6114" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                    <SPLIT distance="100" swimtime="00:01:35.78" />
                    <SPLIT distance="150" swimtime="00:02:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="279" reactiontime="+74" swimtime="00:00:40.01" resultid="3391" heatid="6135" lane="5" entrytime="00:00:33.59" />
                <RESULT eventid="1333" points="356" reactiontime="+92" swimtime="00:00:39.90" resultid="3392" heatid="6206" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1393" points="209" reactiontime="+70" swimtime="00:01:34.68" resultid="3393" heatid="6256" lane="2" entrytime="00:01:18.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="321" reactiontime="+91" swimtime="00:01:32.21" resultid="3394" heatid="6401" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-02" firstname="Konrad" gender="M" lastname="Hasik" nation="POL" athleteid="3395">
              <RESULTS>
                <RESULT eventid="1168" points="698" reactiontime="+85" swimtime="00:01:05.27" resultid="3396" heatid="6095" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="668" reactiontime="+63" swimtime="00:00:29.91" resultid="3397" heatid="6136" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1333" points="665" reactiontime="+81" swimtime="00:00:32.41" resultid="3398" heatid="6215" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1467" points="640" reactiontime="+88" swimtime="00:02:29.77" resultid="3399" heatid="6308" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="150" swimtime="00:01:53.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="558" reactiontime="+83" swimtime="00:00:27.62" resultid="3400" heatid="6356" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1610" points="308" reactiontime="+86" swimtime="00:01:33.54" resultid="3401" heatid="6405" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-05-05" firstname="Robert" gender="M" lastname="Lesiak" nation="POL" athleteid="3402">
              <RESULTS>
                <RESULT eventid="1168" points="375" reactiontime="+92" swimtime="00:01:20.74" resultid="3403" heatid="6094" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="423" reactiontime="+74" swimtime="00:00:34.78" resultid="3404" heatid="6135" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1363" points="427" reactiontime="+93" swimtime="00:00:33.54" resultid="3405" heatid="6234" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1393" points="375" reactiontime="+72" swimtime="00:01:18.54" resultid="3406" heatid="6258" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="3407" heatid="6323" lane="6" entrytime="00:01:14.00" />
                <RESULT eventid="1558" points="587" reactiontime="+63" swimtime="00:02:31.01" resultid="3408" heatid="6381" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:13.58" />
                    <SPLIT distance="150" swimtime="00:01:52.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-08-08" firstname="Damien" gender="M" lastname="Fevier" nation="POL" athleteid="3409">
              <RESULTS>
                <RESULT eventid="1137" points="328" swimtime="00:12:10.43" resultid="3410" heatid="6452" lane="3" entrytime="00:11:27.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                    <SPLIT distance="100" swimtime="00:01:22.18" />
                    <SPLIT distance="200" swimtime="00:02:51.93" />
                    <SPLIT distance="300" swimtime="00:04:24.28" />
                    <SPLIT distance="400" swimtime="00:05:58.78" />
                    <SPLIT distance="500" swimtime="00:07:33.75" />
                    <SPLIT distance="600" swimtime="00:09:08.73" />
                    <SPLIT distance="700" swimtime="00:10:41.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="446" reactiontime="+84" swimtime="00:01:15.78" resultid="3411" heatid="6095" lane="6" entrytime="00:01:11.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="313" reactiontime="+86" swimtime="00:03:05.37" resultid="3412" heatid="6189" lane="2" entrytime="00:02:57.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:21.41" />
                    <SPLIT distance="150" swimtime="00:02:12.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="620" reactiontime="+80" swimtime="00:00:29.74" resultid="3413" heatid="6237" lane="2" entrytime="00:00:29.77" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="3414" heatid="6307" lane="6" entrytime="00:02:47.77" />
                <RESULT eventid="1528" points="540" reactiontime="+82" swimtime="00:00:27.91" resultid="3415" heatid="6359" lane="2" entrytime="00:00:27.27" />
                <RESULT eventid="1610" points="389" reactiontime="+85" swimtime="00:01:26.52" resultid="3416" heatid="6404" lane="6" entrytime="00:01:21.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+57" swimtime="00:01:59.37" resultid="3417" heatid="6525" lane="4" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:03.91" />
                    <SPLIT distance="150" swimtime="00:01:33.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3381" number="1" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3360" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3365" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3347" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1250" swimtime="00:02:09.16" resultid="3419" heatid="6525" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:11.12" />
                    <SPLIT distance="150" swimtime="00:01:41.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3327" number="1" />
                    <RELAYPOSITION athleteid="3335" number="2" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3409" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3376" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+74" swimtime="00:02:15.11" resultid="3421" heatid="6525" lane="6" entrytime="00:02:06.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                    <SPLIT distance="150" swimtime="00:01:44.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3389" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="3343" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="3351" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3395" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+85" swimtime="00:01:48.57" resultid="3418" heatid="6533" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.89" />
                    <SPLIT distance="100" swimtime="00:00:55.59" />
                    <SPLIT distance="150" swimtime="00:01:22.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3395" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="3360" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3365" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3347" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+77" swimtime="00:01:52.65" resultid="3420" heatid="6533" lane="2" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="100" swimtime="00:00:56.96" />
                    <SPLIT distance="150" swimtime="00:01:24.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3327" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3335" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3376" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="3409" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+80" swimtime="00:02:00.00" resultid="3422" heatid="6533" lane="1" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                    <SPLIT distance="100" swimtime="00:00:58.63" />
                    <SPLIT distance="150" swimtime="00:01:27.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3381" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3343" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="3351" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="3402" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ZKSDRZONKÓ" name="ZKS Drzonków" nation="POL" region="LBS">
          <CONTACT city="ŁĘŻYCA" email="piotrbarta@o2.pl" name="BARTA PIOTR" phone="602347348" state="LUBUS" street="ODRZAŃSKA 21" zip="66016" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-18" firstname="PIOTR" gender="M" lastname="BARTA" nation="POL" athleteid="3447">
              <RESULTS>
                <RESULT eventid="1092" points="696" reactiontime="+88" swimtime="00:05:30.94" resultid="3448" heatid="6492" lane="6" entrytime="00:05:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:10.73" />
                    <SPLIT distance="150" swimtime="00:01:57.38" />
                    <SPLIT distance="200" swimtime="00:02:43.17" />
                    <SPLIT distance="250" swimtime="00:03:28.10" />
                    <SPLIT distance="300" swimtime="00:04:14.31" />
                    <SPLIT distance="350" swimtime="00:04:53.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="819" reactiontime="+85" swimtime="00:02:40.68" resultid="3449" heatid="6116" lane="2" entrytime="00:02:48.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:16.61" />
                    <SPLIT distance="150" swimtime="00:01:58.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="690" reactiontime="+80" swimtime="00:00:33.38" resultid="3450" heatid="6215" lane="6" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1467" points="717" reactiontime="+86" swimtime="00:02:32.36" resultid="3451" heatid="6309" lane="6" entrytime="00:02:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:14.45" />
                    <SPLIT distance="150" swimtime="00:01:56.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="790" reactiontime="+74" swimtime="00:01:12.66" resultid="3452" heatid="6407" lane="6" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="643" reactiontime="+90" swimtime="00:04:51.02" resultid="3453" heatid="6568" lane="6" entrytime="00:04:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                    <SPLIT distance="150" swimtime="00:01:43.70" />
                    <SPLIT distance="200" swimtime="00:02:19.92" />
                    <SPLIT distance="250" swimtime="00:02:56.48" />
                    <SPLIT distance="300" swimtime="00:03:33.46" />
                    <SPLIT distance="350" swimtime="00:04:10.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Mielec" nation="POL">
          <CONTACT name="Boicetta" phone="501072284" />
          <ATHLETES>
            <ATHLETE birthdate="1975-05-20" firstname="Sebastian" gender="M" lastname="Boicetta" nation="POL" athleteid="3455">
              <RESULTS>
                <RESULT eventid="1168" points="364" reactiontime="+86" swimtime="00:01:21.74" resultid="3456" heatid="6088" lane="3" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="374" reactiontime="+69" swimtime="00:00:38.13" resultid="3457" heatid="6133" lane="2" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1393" points="359" reactiontime="+67" swimtime="00:01:22.71" resultid="3458" heatid="6254" lane="4" entrytime="00:01:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-22" firstname="Patryk" gender="M" lastname="Małek" nation="POL" athleteid="3459">
              <RESULTS>
                <RESULT eventid="1168" points="477" reactiontime="+78" swimtime="00:01:14.09" resultid="3460" heatid="6092" lane="4" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-4 - przedwczesny start." eventid="1363" reactiontime="+66" status="DSQ" swimtime="00:00:31.19" resultid="3461" heatid="6233" lane="6" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3462" heatid="6357" lane="6" entrytime="00:00:28.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="SiKReT GLIWICE" nation="POL">
          <CONTACT city="GLIWICE" email="j.zagala@ecotrade.pl" internet="www.sikret-plywanie.pl" name="JOANNA ZAGAŁA" phone="601427257" state="ŚLĄSK" street="JAGIELOŃSKA 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="3464">
              <RESULTS>
                <RESULT eventid="1183" points="365" reactiontime="+91" swimtime="00:04:09.62" resultid="3465" heatid="6103" lane="4" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.09" />
                    <SPLIT distance="100" swimtime="00:01:59.59" />
                    <SPLIT distance="150" swimtime="00:03:04.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="462" reactiontime="+91" swimtime="00:00:49.03" resultid="3466" heatid="6196" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1452" points="276" reactiontime="+83" swimtime="00:04:10.36" resultid="3467" heatid="6294" lane="6" entrytime="00:04:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.36" />
                    <SPLIT distance="100" swimtime="00:02:06.14" />
                    <SPLIT distance="150" swimtime="00:03:11.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="231" reactiontime="+85" swimtime="00:01:59.72" resultid="3468" heatid="6313" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="408" reactiontime="+87" swimtime="00:01:52.33" resultid="3469" heatid="6506" lane="5" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="ZAGAŁA" nation="POL" athleteid="3470">
              <RESULTS>
                <RESULT eventid="1153" points="427" reactiontime="+70" swimtime="00:01:40.40" resultid="3471" heatid="6076" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="381" reactiontime="+76" swimtime="00:01:29.70" resultid="3472" heatid="6151" lane="1" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="447" reactiontime="+78" swimtime="00:00:49.57" resultid="3473" heatid="6194" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="1452" points="399" reactiontime="+76" swimtime="00:03:41.46" resultid="3474" heatid="6294" lane="1" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                    <SPLIT distance="100" swimtime="00:01:47.26" />
                    <SPLIT distance="150" swimtime="00:02:49.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="427" reactiontime="+76" swimtime="00:00:38.69" resultid="3475" heatid="6332" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-14" firstname="Danuta" gender="F" lastname="ZIARKO" nation="POL" athleteid="3476">
              <RESULTS>
                <RESULT eventid="1122" points="370" swimtime="00:13:07.45" resultid="3477" heatid="6443" lane="4" entrytime="00:13:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                    <SPLIT distance="100" swimtime="00:01:30.42" />
                    <SPLIT distance="200" swimtime="00:03:07.51" />
                    <SPLIT distance="300" swimtime="00:04:46.95" />
                    <SPLIT distance="400" swimtime="00:06:25.80" />
                    <SPLIT distance="500" swimtime="00:08:03.95" />
                    <SPLIT distance="600" swimtime="00:09:45.80" />
                    <SPLIT distance="700" swimtime="00:11:28.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="265" reactiontime="+99" swimtime="00:03:43.67" resultid="3478" heatid="6182" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.55" />
                    <SPLIT distance="100" swimtime="00:01:41.02" />
                    <SPLIT distance="150" swimtime="00:02:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="449" reactiontime="+89" swimtime="00:00:37.65" resultid="3479" heatid="6221" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1422" points="388" reactiontime="+64" swimtime="00:02:51.65" resultid="3480" heatid="6275" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                    <SPLIT distance="150" swimtime="00:02:07.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="333" reactiontime="+95" swimtime="00:01:32.24" resultid="3481" heatid="6313" lane="3" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="361" reactiontime="+97" swimtime="00:06:16.39" resultid="3482" heatid="6556" lane="2" entrytime="00:06:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                    <SPLIT distance="100" swimtime="00:01:28.23" />
                    <SPLIT distance="150" swimtime="00:02:15.40" />
                    <SPLIT distance="200" swimtime="00:03:03.58" />
                    <SPLIT distance="250" swimtime="00:03:52.83" />
                    <SPLIT distance="300" swimtime="00:04:41.82" />
                    <SPLIT distance="350" swimtime="00:05:30.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Łukasz" gender="M" lastname="STOLARCZYK" nation="POL" athleteid="3483">
              <RESULTS>
                <RESULT eventid="1272" points="697" reactiontime="+79" swimtime="00:00:57.12" resultid="3484" heatid="6178" lane="4" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="746" reactiontime="+75" swimtime="00:00:27.84" resultid="3485" heatid="6239" lane="1" entrytime="00:00:28.05" />
                <RESULT eventid="1498" points="715" reactiontime="+71" swimtime="00:01:02.29" resultid="3486" heatid="6325" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="700" reactiontime="+73" swimtime="00:00:25.98" resultid="3487" heatid="6363" lane="3" entrytime="00:00:25.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-12-05" firstname="Tomasz" gender="M" lastname="PALUCH" nation="POL" athleteid="3488">
              <RESULTS>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="3489" heatid="6178" lane="3" entrytime="00:00:57.00" />
                <RESULT eventid="1528" points="782" reactiontime="+80" swimtime="00:00:25.12" resultid="3490" heatid="6365" lane="2" entrytime="00:00:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-10-06" firstname="Arkadiusz" gender="M" lastname="BEDNAREK" nation="POL" athleteid="3491">
              <RESULTS>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3492" heatid="6204" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1528" points="219" reactiontime="+96" swimtime="00:00:38.38" resultid="3493" heatid="6345" lane="2" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Wojciech" gender="M" lastname="ŁOŻYŃSKI" nation="POL" athleteid="3494">
              <RESULTS>
                <RESULT eventid="1168" points="657" reactiontime="+111" swimtime="00:01:15.35" resultid="3495" heatid="6091" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="3496" heatid="6169" lane="1" entrytime="00:01:07.00" />
                <RESULT eventid="1498" points="608" reactiontime="+91" swimtime="00:01:14.55" resultid="3497" heatid="6321" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-10" firstname="Ioannis" gender="M" lastname="GIOVANIS" nation="POL" athleteid="3498" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+71" swimtime="00:02:10.31" resultid="3502" heatid="6524" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="100" swimtime="00:01:18.09" />
                    <SPLIT distance="150" swimtime="00:01:45.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3494" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3483" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="3491" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="3488" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1415" reactiontime="+97" swimtime="00:02:00.90" resultid="6518" heatid="6530" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                    <SPLIT distance="150" swimtime="00:01:35.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3498" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="3491" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3488" number="3" />
                    <RELAYPOSITION athleteid="3483" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+81" swimtime="00:02:07.09" resultid="3499" heatid="6497" lane="6" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.18" />
                    <SPLIT distance="150" swimtime="00:01:35.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3488" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3470" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="3476" number="3" />
                    <RELAYPOSITION athleteid="3483" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1588" reactiontime="+79" swimtime="00:02:27.28" resultid="3501" heatid="6537" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.87" />
                    <SPLIT distance="100" swimtime="00:01:34.33" />
                    <SPLIT distance="150" swimtime="00:02:02.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3476" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="3464" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3488" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="3483" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Sinnet" nation="POL">
          <CONTACT city="Warszawa" email="piotrbarski@uw.edu.pl" name="Barski" street="Gołkowska 2" />
          <ATHLETES>
            <ATHLETE birthdate="1965-02-17" firstname="Piotr" gender="M" lastname="Barski" nation="POL" athleteid="3504">
              <RESULTS>
                <RESULT eventid="1198" points="816" reactiontime="+86" swimtime="00:02:44.74" resultid="3505" heatid="6114" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:18.30" />
                    <SPLIT distance="150" swimtime="00:02:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="816" reactiontime="+83" swimtime="00:00:58.59" resultid="3506" heatid="6175" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="820" reactiontime="+81" swimtime="00:00:32.82" resultid="3507" heatid="6216" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1363" points="811" reactiontime="+79" swimtime="00:00:29.36" resultid="3508" heatid="6239" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1528" points="794" reactiontime="+76" swimtime="00:00:26.49" resultid="3509" heatid="6362" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1610" points="818" reactiontime="+78" swimtime="00:01:13.51" resultid="3510" heatid="6405" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-25" firstname="Agnieszka" gender="F" lastname="Besler" nation="POL" athleteid="3511">
              <RESULTS>
                <RESULT eventid="1153" points="352" reactiontime="+91" swimtime="00:01:32.03" resultid="3512" heatid="6077" lane="4" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="413" reactiontime="+84" swimtime="00:01:17.95" resultid="3513" heatid="6154" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="440" reactiontime="+80" swimtime="00:00:43.73" resultid="3514" heatid="6198" lane="6" entrytime="00:00:45.70" />
                <RESULT eventid="1595" points="450" reactiontime="+91" swimtime="00:01:33.15" resultid="3515" heatid="6507" lane="4" entrytime="00:01:37.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-18" firstname="Joanna" gender="F" lastname="Janicka" nation="POL" athleteid="3516">
              <RESULTS>
                <RESULT eventid="1257" points="587" reactiontime="+88" swimtime="00:01:08.60" resultid="3517" heatid="6156" lane="2" entrytime="00:01:12.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="648" swimtime="00:00:33.68" resultid="3518" heatid="6223" lane="2" entrytime="00:00:31.25" />
                <RESULT eventid="1513" points="640" reactiontime="+90" swimtime="00:00:30.62" resultid="3519" heatid="6339" lane="4" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STAPOZ" name="Start Poznań" nation="POL" region="WIE">
          <CONTACT city="POZNAŃ" email="ssimasterslukaszewicz@wp.pl" fax="61 8411059" name="ŁUKASZEWICZ PAWEŁ" phone="505186845" state="WIE" street="ZACISZE" street2="2" zip="60-831" />
          <ATHLETES>
            <ATHLETE birthdate="1973-10-22" firstname="Sabina" gender="F" lastname="Rogala-Łukaszewicz" nation="POL" athleteid="3523">
              <RESULTS>
                <RESULT eventid="1153" points="495" reactiontime="+98" swimtime="00:01:25.54" resultid="3524" heatid="6079" lane="2" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="523" reactiontime="+88" swimtime="00:01:11.60" resultid="3525" heatid="6156" lane="4" entrytime="00:01:10.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="486" reactiontime="+90" swimtime="00:00:37.19" resultid="3526" heatid="6220" lane="3" entrytime="00:00:38.16" entrycourse="SCM" />
                <RESULT eventid="1422" points="457" reactiontime="+95" swimtime="00:02:43.26" resultid="3527" heatid="6275" lane="3" entrytime="00:02:51.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:18.31" />
                    <SPLIT distance="150" swimtime="00:02:00.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="561" reactiontime="+82" swimtime="00:00:32.49" resultid="3528" heatid="6338" lane="6" entrytime="00:00:31.96" entrycourse="SCM" />
                <RESULT eventid="1595" points="464" reactiontime="+89" swimtime="00:01:35.77" resultid="3529" heatid="6507" lane="3" entrytime="00:01:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-12-18" firstname="Paweł" gender="M" lastname="Łukaszewicz" nation="POL" athleteid="3530">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="3531" heatid="6088" lane="1" entrytime="00:01:25.00" entrycourse="SCM" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="3532" heatid="6165" lane="5" entrytime="00:01:12.00" entrycourse="SCM" />
                <RESULT eventid="1393" points="531" reactiontime="+68" swimtime="00:01:23.43" resultid="3533" heatid="6254" lane="3" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="467" reactiontime="+101" swimtime="00:02:49.83" resultid="3534" heatid="6283" lane="5" entrytime="00:02:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:01:56.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="533" reactiontime="+73" swimtime="00:03:05.70" resultid="3535" heatid="6376" lane="4" entrytime="00:03:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                    <SPLIT distance="100" swimtime="00:01:29.39" />
                    <SPLIT distance="150" swimtime="00:02:17.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="485" reactiontime="+111" swimtime="00:06:04.16" resultid="3536" heatid="6563" lane="3" entrytime="00:05:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:22.81" />
                    <SPLIT distance="150" swimtime="00:02:09.45" />
                    <SPLIT distance="200" swimtime="00:02:56.70" />
                    <SPLIT distance="250" swimtime="00:03:43.78" />
                    <SPLIT distance="300" swimtime="00:04:31.74" />
                    <SPLIT distance="350" swimtime="00:05:18.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-27" firstname="Krzysztof" gender="M" lastname="Kapałczyński" nation="POL" athleteid="3537">
              <RESULTS>
                <RESULT eventid="1092" points="606" reactiontime="+87" swimtime="00:05:58.92" resultid="3538" heatid="6490" lane="2" entrytime="00:06:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:18.67" />
                    <SPLIT distance="150" swimtime="00:02:05.80" />
                    <SPLIT distance="200" swimtime="00:02:52.98" />
                    <SPLIT distance="250" swimtime="00:03:43.28" />
                    <SPLIT distance="300" swimtime="00:04:34.13" />
                    <SPLIT distance="350" swimtime="00:05:17.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="628" reactiontime="+91" swimtime="00:02:59.81" resultid="3539" heatid="6114" lane="5" entrytime="00:03:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                    <SPLIT distance="100" swimtime="00:01:25.18" />
                    <SPLIT distance="150" swimtime="00:02:13.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="518" reactiontime="+87" swimtime="00:02:56.56" resultid="3540" heatid="6189" lane="1" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:21.95" />
                    <SPLIT distance="150" swimtime="00:02:09.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="582" reactiontime="+86" swimtime="00:02:47.41" resultid="3541" heatid="6306" lane="2" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:18.14" />
                    <SPLIT distance="150" swimtime="00:02:07.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="491" reactiontime="+85" swimtime="00:01:17.75" resultid="3542" heatid="6322" lane="5" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="557" reactiontime="+85" swimtime="00:01:23.52" resultid="3543" heatid="6403" lane="4" entrytime="00:01:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-02" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="3544">
              <RESULTS>
                <RESULT comment="Rekord Polski kat.E" eventid="1092" points="836" reactiontime="+79" swimtime="00:05:22.45" resultid="3545" heatid="6492" lane="1" entrytime="00:05:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:01:55.86" />
                    <SPLIT distance="200" swimtime="00:02:36.82" />
                    <SPLIT distance="250" swimtime="00:03:23.43" />
                    <SPLIT distance="300" swimtime="00:04:10.91" />
                    <SPLIT distance="350" swimtime="00:04:47.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="833" reactiontime="+75" swimtime="00:01:07.59" resultid="3546" heatid="6096" lane="3" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="855" reactiontime="+75" swimtime="00:00:57.69" resultid="3547" heatid="6176" lane="3" entrytime="00:00:58.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="832" reactiontime="+78" swimtime="00:02:10.29" resultid="3548" heatid="6290" lane="2" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:03.16" />
                    <SPLIT distance="150" swimtime="00:01:36.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="763" reactiontime="+77" swimtime="00:00:26.84" resultid="3549" heatid="6361" lane="6" entrytime="00:00:26.70" entrycourse="SCM" />
                <RESULT eventid="1640" points="810" reactiontime="+84" swimtime="00:04:41.89" resultid="3550" heatid="6568" lane="4" entrytime="00:04:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:07.18" />
                    <SPLIT distance="150" swimtime="00:01:42.73" />
                    <SPLIT distance="200" swimtime="00:02:18.89" />
                    <SPLIT distance="250" swimtime="00:02:55.22" />
                    <SPLIT distance="300" swimtime="00:03:31.37" />
                    <SPLIT distance="350" swimtime="00:04:07.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-16" firstname="Wojciech" gender="M" lastname="Dmytrów" nation="POL" athleteid="3551">
              <RESULTS>
                <RESULT eventid="1198" points="674" reactiontime="+83" swimtime="00:03:03.86" resultid="3552" heatid="6112" lane="4" entrytime="00:03:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:01:26.48" />
                    <SPLIT distance="150" swimtime="00:02:14.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="715" reactiontime="+89" swimtime="00:00:36.00" resultid="3553" heatid="6212" lane="6" entrytime="00:00:37.50" entrycourse="SCM" />
                <RESULT eventid="1610" points="773" reactiontime="+76" swimtime="00:01:19.26" resultid="3554" heatid="6402" lane="5" entrytime="00:01:25.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-26" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="3555" />
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="&apos;Start&apos; Wrocław" nation="POL" region="DOL">
          <CONTACT city="WROCŁAW" email="WZSSTART@POST.PL" fax="071 34 372 81" internet="www.start.wroclaw.pl" name="&apos;START&apos; WROCŁAW" phone="071 34 302 31" state="DOL" street="NOTECKA 12" zip="54-128" />
          <ATHLETES>
            <ATHLETE birthdate="1974-04-30" firstname="Sebastian" gender="M" lastname="Szymański" nation="POL" athleteid="3557">
              <RESULTS>
                <RESULT eventid="1228" points="521" reactiontime="+78" swimtime="00:00:34.14" resultid="3558" heatid="6134" lane="2" entrytime="00:00:34.34" entrycourse="SCM" />
                <RESULT eventid="1272" points="588" reactiontime="+92" swimtime="00:01:01.36" resultid="3559" heatid="6172" lane="4" entrytime="00:01:02.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="586" reactiontime="+99" swimtime="00:00:30.04" resultid="3560" heatid="6234" lane="4" entrytime="00:00:30.78" entrycourse="SCM" />
                <RESULT eventid="1393" points="459" reactiontime="+105" swimtime="00:01:16.20" resultid="3561" heatid="6258" lane="2" entrytime="00:01:14.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="576" reactiontime="+97" swimtime="00:01:08.60" resultid="3562" heatid="6323" lane="1" entrytime="00:01:12.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="562" reactiontime="+98" swimtime="00:00:28.04" resultid="3563" heatid="6356" lane="1" entrytime="00:00:28.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-08-29" firstname="Bartosz" gender="M" lastname="Bogucki" nation="POL" athleteid="3564">
              <RESULTS>
                <RESULT eventid="1363" points="469" reactiontime="+66" swimtime="00:00:32.50" resultid="3565" heatid="6232" lane="3" entrytime="00:00:31.31" entrycourse="SCM" />
                <RESULT eventid="1393" points="367" reactiontime="+66" swimtime="00:01:19.10" resultid="3566" heatid="6257" lane="2" entrytime="00:01:16.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="495" reactiontime="+81" swimtime="00:00:29.15" resultid="3567" heatid="6355" lane="4" entrytime="00:00:28.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Toruńczyk Masters Toruń" nation="POL" region="KUJ">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1952-07-06" firstname="Andrzej" gender="M" lastname="Szufarski" nation="POL" athleteid="3569">
              <RESULTS>
                <RESULT eventid="1198" points="443" reactiontime="+111" swimtime="00:03:51.51" resultid="3570" heatid="6110" lane="3" entrytime="00:03:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.65" />
                    <SPLIT distance="100" swimtime="00:01:47.19" />
                    <SPLIT distance="150" swimtime="00:02:48.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="404" reactiontime="+102" swimtime="00:00:46.34" resultid="3571" heatid="6206" lane="5" entrytime="00:00:44.50" />
                <RESULT eventid="1393" points="274" reactiontime="+105" swimtime="00:01:53.20" resultid="3572" heatid="6252" lane="5" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="3573" heatid="6318" lane="1" entrytime="00:01:38.50" />
                <RESULT eventid="1610" status="DNS" swimtime="00:00:00.00" resultid="3574" heatid="6398" lane="6" entrytime="00:01:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-03" firstname="Artur" gender="M" lastname="Kłosiński" nation="POL" athleteid="3575">
              <RESULTS>
                <RESULT eventid="1228" points="473" reactiontime="+61" swimtime="00:00:33.51" resultid="3576" heatid="6131" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1272" points="569" reactiontime="+81" swimtime="00:01:01.11" resultid="3577" heatid="6176" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="566" reactiontime="+82" swimtime="00:00:35.61" resultid="3578" heatid="6213" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1393" status="DNS" swimtime="00:00:00.00" resultid="3579" heatid="6259" lane="2" entrytime="00:01:11.00" />
                <RESULT eventid="1528" points="612" reactiontime="+80" swimtime="00:00:27.16" resultid="3580" heatid="6363" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1610" points="490" reactiontime="+82" swimtime="00:01:22.28" resultid="3581" heatid="6405" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="3582">
              <RESULTS>
                <RESULT eventid="1168" points="621" reactiontime="+82" swimtime="00:01:24.26" resultid="3583" heatid="6089" lane="5" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="581" reactiontime="+79" swimtime="00:01:14.73" resultid="3584" heatid="6164" lane="5" entrytime="00:01:13.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="668" reactiontime="+50" swimtime="00:00:34.73" resultid="3585" heatid="6229" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1498" points="427" reactiontime="+74" swimtime="00:01:33.03" resultid="3586" heatid="6319" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="608" reactiontime="+76" swimtime="00:00:32.21" resultid="3587" heatid="6349" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1467" points="524" reactiontime="+88" swimtime="00:03:19.76" resultid="6023" heatid="6303" lane="1" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                    <SPLIT distance="100" swimtime="00:01:37.54" />
                    <SPLIT distance="150" swimtime="00:02:34.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="3596">
              <RESULTS>
                <RESULT eventid="1228" points="277" reactiontime="+80" swimtime="00:00:58.58" resultid="3597" heatid="6127" lane="5" entrytime="00:00:56.52" />
                <RESULT eventid="1272" points="325" reactiontime="+121" swimtime="00:01:37.52" resultid="3598" heatid="6160" lane="5" entrytime="00:01:34.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="232" reactiontime="+70" swimtime="00:02:17.46" resultid="3599" heatid="6250" lane="3" entrytime="00:02:08.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="246" reactiontime="+110" swimtime="00:04:06.79" resultid="3600" heatid="6278" lane="3" entrytime="00:03:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.72" />
                    <SPLIT distance="100" swimtime="00:01:58.13" />
                    <SPLIT distance="150" swimtime="00:03:03.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="433" reactiontime="+122" swimtime="00:00:39.84" resultid="3601" heatid="6342" lane="5" entrytime="00:00:59.65" />
                <RESULT eventid="1558" points="248" reactiontime="+86" swimtime="00:04:54.94" resultid="3602" heatid="6373" lane="6" entrytime="00:04:35.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.47" />
                    <SPLIT distance="100" swimtime="00:02:24.82" />
                    <SPLIT distance="150" swimtime="00:03:42.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-23" firstname="Marcin" gender="M" lastname="Mykowski" nation="POL" athleteid="3603">
              <RESULTS>
                <RESULT eventid="1228" points="667" reactiontime="+61" swimtime="00:00:29.87" resultid="3604" heatid="6137" lane="6" entrytime="00:00:31.50" />
                <RESULT eventid="1272" points="694" reactiontime="+77" swimtime="00:00:57.19" resultid="3605" heatid="6177" lane="2" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="636" swimtime="00:01:05.89" resultid="3606" heatid="6261" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="3607" heatid="6291" lane="1" entrytime="00:02:10.00" />
                <RESULT eventid="1558" points="648" reactiontime="+70" swimtime="00:02:26.04" resultid="3608" heatid="6380" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:12.28" />
                    <SPLIT distance="150" swimtime="00:01:49.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-27" firstname="Magdalena" gender="F" lastname="Rogozińska" nation="POL" athleteid="3609">
              <RESULTS>
                <RESULT eventid="1153" points="528" reactiontime="+92" swimtime="00:01:23.76" resultid="3610" heatid="6080" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="458" reactiontime="+94" swimtime="00:03:28.00" resultid="3611" heatid="6106" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                    <SPLIT distance="100" swimtime="00:01:40.52" />
                    <SPLIT distance="150" swimtime="00:02:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="477" reactiontime="+93" swimtime="00:00:42.81" resultid="3612" heatid="6200" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1452" points="464" reactiontime="+115" swimtime="00:03:03.51" resultid="3613" heatid="6295" lane="2" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:28.59" />
                    <SPLIT distance="150" swimtime="00:02:22.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="477" reactiontime="+91" swimtime="00:00:34.30" resultid="3614" heatid="6337" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1595" points="495" reactiontime="+97" swimtime="00:01:33.76" resultid="3615" heatid="6508" lane="3" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-27" firstname="Mariola" gender="F" lastname="Kutc" nation="POL" athleteid="3616">
              <RESULTS>
                <RESULT eventid="1153" points="476" reactiontime="+109" swimtime="00:01:36.81" resultid="3617" heatid="6077" lane="3" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="459" reactiontime="+94" swimtime="00:00:44.85" resultid="3618" heatid="6122" lane="1" entrytime="00:00:44.00" />
                <RESULT eventid="1348" points="517" swimtime="00:00:41.07" resultid="3619" heatid="6220" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1378" points="440" reactiontime="+86" swimtime="00:01:41.53" resultid="3620" heatid="6245" lane="2" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="462" reactiontime="+120" swimtime="00:01:35.08" resultid="3621" heatid="6314" lane="6" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="3622" heatid="6507" lane="1" entrytime="00:01:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-16" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="3623">
              <RESULTS>
                <RESULT eventid="1122" points="360" swimtime="00:12:17.54" resultid="3624" heatid="6445" lane="6" entrytime="00:11:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                    <SPLIT distance="100" swimtime="00:01:23.81" />
                    <SPLIT distance="150" swimtime="00:02:08.37" />
                    <SPLIT distance="200" swimtime="00:02:53.90" />
                    <SPLIT distance="250" swimtime="00:03:39.44" />
                    <SPLIT distance="300" swimtime="00:04:24.88" />
                    <SPLIT distance="350" swimtime="00:05:10.96" />
                    <SPLIT distance="400" swimtime="00:05:57.28" />
                    <SPLIT distance="450" swimtime="00:06:44.80" />
                    <SPLIT distance="500" swimtime="00:07:31.92" />
                    <SPLIT distance="550" swimtime="00:08:19.65" />
                    <SPLIT distance="600" swimtime="00:09:07.52" />
                    <SPLIT distance="650" swimtime="00:09:55.77" />
                    <SPLIT distance="700" swimtime="00:10:43.46" />
                    <SPLIT distance="750" swimtime="00:11:32.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="524" reactiontime="+80" swimtime="00:01:23.06" resultid="3625" heatid="6080" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="480" reactiontime="+73" swimtime="00:01:11.27" resultid="3626" heatid="6158" lane="1" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - przedwczesny start." eventid="1422" reactiontime="+56" status="DSQ" swimtime="00:02:45.85" resultid="3627" heatid="6276" lane="4" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:15.68" />
                    <SPLIT distance="150" swimtime="00:01:59.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="415" reactiontime="+72" swimtime="00:03:06.21" resultid="3628" heatid="6297" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                    <SPLIT distance="150" swimtime="00:02:20.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="373" reactiontime="+75" swimtime="00:03:08.40" resultid="3629" heatid="6371" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                    <SPLIT distance="100" swimtime="00:01:33.31" />
                    <SPLIT distance="150" swimtime="00:02:21.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="400" reactiontime="+75" swimtime="00:05:44.14" resultid="3630" heatid="6557" lane="3" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:20.43" />
                    <SPLIT distance="150" swimtime="00:02:04.07" />
                    <SPLIT distance="200" swimtime="00:02:48.49" />
                    <SPLIT distance="250" swimtime="00:03:32.47" />
                    <SPLIT distance="300" swimtime="00:04:17.03" />
                    <SPLIT distance="350" swimtime="00:05:01.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-14" firstname="Marta" gender="F" lastname="Lord" nation="POL" athleteid="3631">
              <RESULTS>
                <RESULT eventid="1153" points="598" reactiontime="+87" swimtime="00:01:17.16" resultid="3632" heatid="6080" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="627" reactiontime="+90" swimtime="00:00:35.62" resultid="3633" heatid="6124" lane="2" entrytime="00:00:36.68" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="3634" heatid="6200" lane="2" entrytime="00:00:40.30" />
                <RESULT eventid="1378" points="624" reactiontime="+85" swimtime="00:01:16.69" resultid="3635" heatid="6247" lane="3" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. B" eventid="1543" points="659" reactiontime="+94" swimtime="00:02:39.84" resultid="3636" heatid="6371" lane="6" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                    <SPLIT distance="100" swimtime="00:01:18.66" />
                    <SPLIT distance="150" swimtime="00:02:00.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-04" firstname="Karol" gender="M" lastname="Twarowski" nation="POL" athleteid="3637">
              <RESULTS>
                <RESULT eventid="1137" points="690" swimtime="00:09:24.06" resultid="3638" heatid="6455" lane="4" entrytime="00:10:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:01.71" />
                    <SPLIT distance="200" swimtime="00:02:11.10" />
                    <SPLIT distance="300" swimtime="00:03:20.70" />
                    <SPLIT distance="400" swimtime="00:04:31.24" />
                    <SPLIT distance="500" swimtime="00:05:42.36" />
                    <SPLIT distance="600" swimtime="00:06:54.92" />
                    <SPLIT distance="700" swimtime="00:08:08.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="760" reactiontime="+82" swimtime="00:01:03.85" resultid="3639" heatid="6097" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="754" reactiontime="+77" swimtime="00:00:55.64" resultid="3640" heatid="6177" lane="4" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="682" reactiontime="+78" swimtime="00:01:04.36" resultid="3641" heatid="6260" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="756" reactiontime="+85" swimtime="00:02:02.56" resultid="3642" heatid="6290" lane="1" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="100" swimtime="00:00:59.01" />
                    <SPLIT distance="150" swimtime="00:01:30.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="684" reactiontime="+83" swimtime="00:01:03.23" resultid="3643" heatid="6323" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="732" reactiontime="+83" swimtime="00:02:20.26" resultid="3644" heatid="6381" lane="2" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="100" swimtime="00:01:07.03" />
                    <SPLIT distance="150" swimtime="00:01:42.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="3645">
              <RESULTS>
                <RESULT eventid="1302" points="353" reactiontime="+88" swimtime="00:02:57.94" resultid="3646" heatid="6188" lane="5" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                    <SPLIT distance="100" swimtime="00:01:20.32" />
                    <SPLIT distance="150" swimtime="00:02:08.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="484" reactiontime="+82" swimtime="00:00:32.17" resultid="3647" heatid="6231" lane="4" entrytime="00:00:32.50" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="3648" heatid="6284" lane="2" entrytime="00:02:35.00" />
                <RESULT eventid="1498" points="439" reactiontime="+81" swimtime="00:01:13.30" resultid="3649" heatid="6322" lane="4" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="353" reactiontime="+83" swimtime="00:05:40.31" resultid="3650" heatid="6565" lane="2" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="100" swimtime="00:01:19.66" />
                    <SPLIT distance="150" swimtime="00:02:03.95" />
                    <SPLIT distance="200" swimtime="00:02:47.95" />
                    <SPLIT distance="250" swimtime="00:03:31.70" />
                    <SPLIT distance="300" swimtime="00:04:14.49" />
                    <SPLIT distance="350" swimtime="00:04:57.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-10-22" firstname="Magdalena" gender="F" lastname="Bolewska" nation="POL" athleteid="3651">
              <RESULTS>
                <RESULT eventid="1183" points="680" reactiontime="+94" swimtime="00:02:59.44" resultid="3652" heatid="6107" lane="2" entrytime="00:02:55.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:01:25.97" />
                    <SPLIT distance="150" swimtime="00:02:12.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="639" reactiontime="+89" swimtime="00:01:06.70" resultid="3653" heatid="6157" lane="2" entrytime="00:01:07.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="737" reactiontime="+86" swimtime="00:00:37.73" resultid="3654" heatid="6201" lane="6" entrytime="00:00:37.56" />
                <RESULT eventid="1452" points="635" reactiontime="+90" swimtime="00:02:45.11" resultid="3655" heatid="6298" lane="6" entrytime="00:02:48.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:03.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="578" reactiontime="+89" swimtime="00:01:15.79" resultid="3656" heatid="6315" lane="2" entrytime="00:01:14.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="645" reactiontime="+85" swimtime="00:01:21.83" resultid="3657" heatid="6510" lane="2" entrytime="00:01:21.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-16" firstname="Maciej" gender="M" lastname="Kujawa" nation="POL" athleteid="3658">
              <RESULTS>
                <RESULT eventid="1168" points="608" reactiontime="+104" swimtime="00:01:20.25" resultid="3659" heatid="6091" lane="5" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="606" reactiontime="+99" swimtime="00:00:39.24" resultid="3660" heatid="6209" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1610" points="610" reactiontime="+103" swimtime="00:01:27.58" resultid="3661" heatid="6400" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="6540">
              <RESULTS>
                <RESULT eventid="1302" points="156" reactiontime="+117" swimtime="00:05:00.72" resultid="6541" heatid="6184" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.02" />
                    <SPLIT distance="100" swimtime="00:02:25.82" />
                    <SPLIT distance="150" swimtime="00:03:45.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="120" reactiontime="+83" swimtime="00:02:29.01" resultid="6542" heatid="6250" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="225" swimtime="00:03:52.15" resultid="6543" heatid="6279" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                    <SPLIT distance="100" swimtime="00:01:51.21" />
                    <SPLIT distance="150" swimtime="00:02:53.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="132" reactiontime="+92" swimtime="00:05:17.66" resultid="6544" heatid="6372" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.81" />
                    <SPLIT distance="100" swimtime="00:02:36.21" />
                    <SPLIT distance="150" swimtime="00:03:58.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" status="DNS" swimtime="00:00:00.00" resultid="6545" heatid="6559" lane="4" />
                <RESULT eventid="1228" points="120" reactiontime="+103" swimtime="00:01:07.74" resultid="6548" heatid="6126" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+67" swimtime="00:02:04.04" resultid="3664" heatid="6524" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:06.56" />
                    <SPLIT distance="150" swimtime="00:01:38.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3603" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3575" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="3645" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="3637" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1415" reactiontime="+80" swimtime="00:01:47.75" resultid="3665" heatid="6534" lane="6" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                    <SPLIT distance="100" swimtime="00:00:52.17" />
                    <SPLIT distance="150" swimtime="00:01:21.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3575" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3645" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="3603" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3637" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+83" swimtime="00:02:42.08" resultid="3666" heatid="6522" lane="1" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                    <SPLIT distance="100" swimtime="00:01:28.35" />
                    <SPLIT distance="150" swimtime="00:02:03.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3658" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="3569" number="2" reactiontime="+97" />
                    <RELAYPOSITION athleteid="3582" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="3596" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1415" reactiontime="+100" swimtime="00:02:24.44" resultid="3667" heatid="6531" lane="6" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:53.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3569" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="3596" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="3658" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="3582" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1408" reactiontime="+83" swimtime="00:02:13.50" resultid="3662" heatid="6528" lane="5" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                    <SPLIT distance="100" swimtime="00:01:04.23" />
                    <SPLIT distance="150" swimtime="00:01:43.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3651" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="3631" number="2" reactiontime="+89" />
                    <RELAYPOSITION athleteid="3609" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3616" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1243" reactiontime="+94" swimtime="00:02:33.37" resultid="3663" heatid="6520" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.50" />
                    <SPLIT distance="100" swimtime="00:01:27.67" />
                    <SPLIT distance="150" swimtime="00:02:03.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3616" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="3609" number="2" reactiontime="+94" />
                    <RELAYPOSITION athleteid="3631" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="3651" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+88" swimtime="00:02:05.96" resultid="3668" heatid="6538" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:39.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3603" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="3631" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="3651" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3637" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="T.P.Masters Opole" nation="POL">
          <CONTACT city="OPOLE" email="opolbud@onet.eu" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1931-01-01" firstname="JÓZEF" gender="M" lastname="KASPEREK" nation="POL" athleteid="3692">
              <RESULTS>
                <RESULT eventid="1393" points="145" reactiontime="+56" swimtime="00:02:56.58" resultid="3693" heatid="6250" lane="2" entrytime="00:03:03.00" />
                <RESULT eventid="1437" points="120" reactiontime="+112" swimtime="00:06:30.06" resultid="3694" heatid="6278" lane="5" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.35" />
                    <SPLIT distance="100" swimtime="00:03:05.50" />
                    <SPLIT distance="150" swimtime="00:04:53.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="TADEUSZ" gender="M" lastname="WITKOWSKI" nation="POL" athleteid="3695">
              <RESULTS>
                <RESULT eventid="1092" points="329" reactiontime="+132" swimtime="00:09:57.42" resultid="3696" heatid="6485" lane="5" entrytime="00:09:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.93" />
                    <SPLIT distance="100" swimtime="00:02:34.50" />
                    <SPLIT distance="150" swimtime="00:03:52.04" />
                    <SPLIT distance="200" swimtime="00:06:33.37" />
                    <SPLIT distance="250" swimtime="00:09:00.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="549" reactiontime="+161" swimtime="00:00:48.26" resultid="3697" heatid="6128" lane="4" entrytime="00:00:49.00" />
                <RESULT eventid="1272" points="543" reactiontime="+115" swimtime="00:01:30.72" resultid="3698" heatid="6161" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="471" reactiontime="+117" swimtime="00:00:51.50" resultid="3699" heatid="6204" lane="3" entrytime="00:00:49.50" />
                <RESULT comment="Rekord Polski kat. K" eventid="1393" points="527" reactiontime="+88" swimtime="00:01:49.02" resultid="3700" heatid="6251" lane="3" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="792" reactiontime="+101" swimtime="00:00:35.43" resultid="3701" heatid="6345" lane="4" entrytime="00:00:35.00" />
                <RESULT comment="Rekord Polski kat. K" eventid="1558" points="506" reactiontime="+91" swimtime="00:03:55.63" resultid="3702" heatid="6373" lane="5" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:56.60" />
                    <SPLIT distance="100" swimtime="00:02:58.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="ROMAN" gender="M" lastname="BIRECKI" nation="POL" athleteid="3703">
              <RESULTS>
                <RESULT eventid="1168" points="545" reactiontime="+103" swimtime="00:01:23.24" resultid="3704" heatid="6088" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. G" eventid="1302" points="567" reactiontime="+94" swimtime="00:03:03.92" resultid="3705" heatid="6188" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:01:26.42" />
                    <SPLIT distance="150" swimtime="00:02:15.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="497" reactiontime="+98" swimtime="00:00:35.43" resultid="3706" heatid="6227" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1437" points="563" reactiontime="+104" swimtime="00:02:39.57" resultid="3707" heatid="6282" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:17.01" />
                    <SPLIT distance="150" swimtime="00:02:00.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="JANUSZ" gender="M" lastname="GARBARCZUK" nation="POL" athleteid="3708">
              <RESULTS>
                <RESULT eventid="1228" points="355" reactiontime="+90" swimtime="00:00:47.20" resultid="3709" heatid="6129" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1393" points="304" reactiontime="+81" swimtime="00:01:49.44" resultid="3710" heatid="6252" lane="2" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="MIROSŁAW" gender="M" lastname="URBANIAK" nation="POL" athleteid="3711">
              <RESULTS>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="3712" heatid="6160" lane="1" entrytime="00:01:50.00" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3713" heatid="6206" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="MAREK" gender="M" lastname="CHMIEL" nation="POL" athleteid="3714">
              <RESULTS>
                <RESULT eventid="1333" points="372" swimtime="00:00:42.69" resultid="3715" heatid="6208" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1528" points="353" reactiontime="+96" swimtime="00:00:34.69" resultid="3716" heatid="6346" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="OLGIERD" gender="M" lastname="MIKOSZA" nation="POL" athleteid="3717">
              <RESULTS>
                <RESULT eventid="1228" points="634" reactiontime="+76" swimtime="00:00:38.91" resultid="3718" heatid="6132" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1272" points="663" reactiontime="+50" swimtime="00:01:11.51" resultid="3719" heatid="6168" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="605" reactiontime="+76" swimtime="00:01:26.98" resultid="3720" heatid="6255" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="556" reactiontime="+92" swimtime="00:02:51.69" resultid="3721" heatid="6282" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="150" swimtime="00:02:05.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="729" reactiontime="+87" swimtime="00:00:30.31" resultid="3722" heatid="6352" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1558" points="564" reactiontime="+87" swimtime="00:03:15.90" resultid="3723" heatid="6376" lane="1" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.47" />
                    <SPLIT distance="100" swimtime="00:01:35.47" />
                    <SPLIT distance="150" swimtime="00:02:28.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="OSKAR" gender="M" lastname="ORSKI" nation="POL" athleteid="3724">
              <RESULTS>
                <RESULT eventid="1272" points="481" reactiontime="+100" swimtime="00:01:09.89" resultid="3725" heatid="6166" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="ZBIGNIEW" gender="M" lastname="JANUSZKIEWICZ" nation="POL" athleteid="3726">
              <RESULTS>
                <RESULT eventid="1228" points="898" reactiontime="+61" swimtime="00:00:31.73" resultid="3727" heatid="6136" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1393" points="937" reactiontime="+67" swimtime="00:01:08.65" resultid="3728" heatid="6259" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="938" reactiontime="+67" swimtime="00:02:32.15" resultid="3729" heatid="6380" lane="2" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:13.50" />
                    <SPLIT distance="150" swimtime="00:01:53.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="ZBIGNIEW" gender="M" lastname="KRASNODĘBSKI" nation="POL" athleteid="3730">
              <RESULTS>
                <RESULT eventid="1333" points="537" reactiontime="+96" swimtime="00:00:40.85" resultid="3731" heatid="6210" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1610" points="536" reactiontime="+103" swimtime="00:01:31.45" resultid="3732" heatid="6401" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="JERZY" gender="M" lastname="MINKIEWICZ" nation="POL" athleteid="3733">
              <RESULTS>
                <RESULT eventid="1168" points="528" reactiontime="+84" swimtime="00:01:24.13" resultid="3734" heatid="6088" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="618" reactiontime="+87" swimtime="00:01:08.87" resultid="3735" heatid="6168" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="492" reactiontime="+90" swimtime="00:00:35.56" resultid="3736" heatid="6229" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1393" points="421" reactiontime="+76" swimtime="00:01:30.14" resultid="3737" heatid="6254" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="352" reactiontime="+100" swimtime="00:01:31.10" resultid="3738" heatid="6319" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="453" reactiontime="+78" swimtime="00:03:15.98" resultid="3739" heatid="6375" lane="2" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.39" />
                    <SPLIT distance="100" swimtime="00:01:38.11" />
                    <SPLIT distance="150" swimtime="00:02:28.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+62" swimtime="00:02:16.68" resultid="3740" heatid="6523" lane="3" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:11.94" />
                    <SPLIT distance="150" swimtime="00:01:47.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3726" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="3730" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3703" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3724" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1415" reactiontime="+91" swimtime="00:02:01.43" resultid="3741" heatid="6532" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:04.99" />
                    <SPLIT distance="150" swimtime="00:01:34.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3726" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="3703" number="2" reactiontime="+86" />
                    <RELAYPOSITION athleteid="3724" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3717" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+67" swimtime="00:02:41.85" resultid="3742" heatid="6522" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                    <SPLIT distance="100" swimtime="00:01:27.70" />
                    <SPLIT distance="150" swimtime="00:02:04.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3717" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3708" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3733" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="3695" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1415" swimtime="00:02:21.16" resultid="3743" heatid="6531" lane="2" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="100" swimtime="00:01:15.21" />
                    <SPLIT distance="150" swimtime="00:01:49.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3695" number="1" />
                    <RELAYPOSITION athleteid="3708" number="2" />
                    <RELAYPOSITION athleteid="3730" number="3" />
                    <RELAYPOSITION athleteid="3733" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="TS Wisła Kraków" nation="POL">
          <CONTACT name="aa" />
          <ATHLETES>
            <ATHLETE birthdate="1930-01-01" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="3760">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. L" eventid="1092" points="1292" reactiontime="+119" swimtime="00:08:22.06" resultid="3761" heatid="6485" lane="2" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.78" />
                    <SPLIT distance="100" swimtime="00:02:04.44" />
                    <SPLIT distance="150" swimtime="00:03:05.36" />
                    <SPLIT distance="200" swimtime="00:04:08.46" />
                    <SPLIT distance="250" swimtime="00:05:20.78" />
                    <SPLIT distance="300" swimtime="00:06:31.23" />
                    <SPLIT distance="350" swimtime="00:07:25.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="897" reactiontime="+105" swimtime="00:01:44.53" resultid="3762" heatid="6085" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="683" reactiontime="+113" swimtime="00:01:27.84" resultid="3763" heatid="6160" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="551" reactiontime="+109" swimtime="00:00:53.88" resultid="3764" heatid="6225" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1437" points="838" swimtime="00:03:24.21" resultid="3765" heatid="6283" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                    <SPLIT distance="100" swimtime="00:01:37.36" />
                    <SPLIT distance="150" swimtime="00:02:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="669" reactiontime="+109" swimtime="00:00:37.90" resultid="3766" heatid="6344" lane="6" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Janusz" gender="M" lastname="Konstanty" nation="POL" athleteid="3767">
              <RESULTS>
                <RESULT eventid="1168" points="632" reactiontime="+89" swimtime="00:01:19.26" resultid="3768" heatid="6090" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="707" reactiontime="+73" swimtime="00:00:35.82" resultid="3769" heatid="6132" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1393" points="653" reactiontime="+83" swimtime="00:01:17.85" resultid="3770" heatid="6256" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="676" reactiontime="+94" swimtime="00:02:56.28" resultid="3771" heatid="6304" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:20.95" />
                    <SPLIT distance="150" swimtime="00:02:14.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="654" reactiontime="+80" swimtime="00:02:53.49" resultid="3772" heatid="6377" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                    <SPLIT distance="100" swimtime="00:01:23.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Paweł" gender="M" lastname="Lesiakowski" nation="POL" athleteid="3773">
              <RESULTS>
                <RESULT eventid="1333" points="612" reactiontime="+81" swimtime="00:00:40.34" resultid="3774" heatid="6207" lane="3" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="3775">
              <RESULTS>
                <RESULT eventid="1058" points="600" reactiontime="+91" swimtime="00:06:54.81" resultid="3776" heatid="6428" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                    <SPLIT distance="100" swimtime="00:01:33.97" />
                    <SPLIT distance="150" swimtime="00:02:27.48" />
                    <SPLIT distance="200" swimtime="00:03:20.16" />
                    <SPLIT distance="250" swimtime="00:04:20.76" />
                    <SPLIT distance="300" swimtime="00:05:22.40" />
                    <SPLIT distance="350" swimtime="00:06:08.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="645" reactiontime="+104" swimtime="00:01:27.47" resultid="3777" heatid="6074" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="549" reactiontime="+108" swimtime="00:03:29.55" resultid="3778" heatid="6181" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                    <SPLIT distance="100" swimtime="00:01:37.10" />
                    <SPLIT distance="150" swimtime="00:02:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="568" reactiontime="+103" swimtime="00:00:39.81" resultid="3779" heatid="6218" lane="6" />
                <RESULT eventid="1452" points="583" reactiontime="+106" swimtime="00:03:15.20" resultid="3780" heatid="6293" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:01:32.19" />
                    <SPLIT distance="150" swimtime="00:02:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="523" reactiontime="+87" swimtime="00:01:31.24" resultid="3781" heatid="6312" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - przedwczesny start." eventid="1513" reactiontime="+98" status="DSQ" swimtime="00:00:34.96" resultid="3782" heatid="6328" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04514" name="Uks 307" nation="POL" region="MAZ">
          <CONTACT name="Ilczyszyn" />
          <ATHLETES>
            <ATHLETE birthdate="1983-07-13" firstname="Krzysztof" gender="M" lastname="Ilczyszyn" nation="POL" athleteid="3784">
              <RESULTS>
                <RESULT eventid="1168" points="465" reactiontime="+83" swimtime="00:01:14.74" resultid="3785" heatid="6092" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="526" reactiontime="+44" swimtime="00:01:02.63" resultid="3786" heatid="6171" lane="2" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="573" reactiontime="+78" swimtime="00:00:30.53" resultid="3787" heatid="6235" lane="5" entrytime="00:00:30.20" />
                <RESULT eventid="1437" points="419" reactiontime="+81" swimtime="00:02:27.86" resultid="3788" heatid="6285" lane="4" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:11.19" />
                    <SPLIT distance="150" swimtime="00:01:50.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="3789" heatid="6321" lane="3" entrytime="00:01:16.00" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3790" heatid="6359" lane="1" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZS SUM" name="AZS Śląski Uniwersytet Medyczny" nation="POL" region="SLA" shortname="AZS Śląski Uniwersytet Medyczn">
          <CONTACT city="Chorzów" email="karol.palka@gmail.com" name="Karol Pałka" phone="693815255" state="ŚLĄSK" street="Śląska 7/1" zip="41-500" />
          <ATHLETES>
            <ATHLETE birthdate="1990-03-18" firstname="Karol" gender="M" lastname="Pałka" nation="POL" athleteid="3792">
              <RESULTS>
                <RESULT eventid="1198" points="417" reactiontime="+85" swimtime="00:03:00.36" resultid="3793" heatid="6116" lane="5" entrytime="00:02:48.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                    <SPLIT distance="100" swimtime="00:01:23.43" />
                    <SPLIT distance="150" swimtime="00:02:11.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="524" reactiontime="+80" swimtime="00:00:35.12" resultid="3794" heatid="6216" lane="1" entrytime="00:00:32.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-10" firstname="Anna" gender="F" lastname="Szczegielniak" nation="POL" athleteid="3795">
              <RESULTS>
                <RESULT eventid="1318" points="185" reactiontime="+131" swimtime="00:00:57.53" resultid="3796" heatid="6197" lane="5" entrytime="00:00:49.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SOPMAST" name="Sopot Masters" nation="POL" region="POM">
          <CONTACT city="SOPOT" email="sopotmasters@o2.pl" internet="www.sopotmasters.pl" name="Gorbaczow Mirosław" phone="696 258 185" state="POMOR" street="ul. Haffnera 57" zip="81-715" />
          <ATHLETES>
            <ATHLETE birthdate="1964-08-04" firstname="JOANNA" gender="F" lastname="PUCHALSKA" nation="POL" athleteid="3798">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. E" eventid="1058" points="1017" reactiontime="+88" swimtime="00:05:41.67" resultid="3799" heatid="6431" lane="3" entrytime="00:05:47.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                    <SPLIT distance="150" swimtime="00:02:00.49" />
                    <SPLIT distance="200" swimtime="00:02:46.04" />
                    <SPLIT distance="250" swimtime="00:03:33.88" />
                    <SPLIT distance="300" swimtime="00:04:22.36" />
                    <SPLIT distance="350" swimtime="00:05:02.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="1000" reactiontime="+97" swimtime="00:02:43.80" resultid="3801" heatid="6182" lane="3" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:17.32" />
                    <SPLIT distance="150" swimtime="00:01:59.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="678" swimtime="00:00:34.71" resultid="3802" heatid="6222" lane="2" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1452" status="DNS" swimtime="00:00:00.00" resultid="3803" heatid="6298" lane="2" entrytime="00:02:45.00" entrycourse="SCM" />
                <RESULT eventid="1483" status="DNS" swimtime="00:00:00.00" resultid="3804" heatid="6315" lane="4" entrytime="00:01:14.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-12-28" firstname="DARIUSZ" gender="M" lastname="GORBACZOW" nation="POL" athleteid="3806">
              <RESULTS>
                <RESULT eventid="1228" points="819" reactiontime="+92" swimtime="00:00:32.72" resultid="3807" heatid="6134" lane="1" entrytime="00:00:34.50" entrycourse="SCM" />
                <RESULT eventid="1363" points="747" reactiontime="+47" swimtime="00:00:30.55" resultid="3808" heatid="6233" lane="2" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1393" points="631" reactiontime="+84" swimtime="00:01:18.31" resultid="3809" heatid="6257" lane="3" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="702" reactiontime="+83" swimtime="00:00:28.54" resultid="3810" heatid="6355" lane="1" entrytime="00:00:28.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-10-13" firstname="MIROSŁAW" gender="M" lastname="GORBACZOW" nation="POL" athleteid="3811">
              <RESULTS>
                <RESULT eventid="1092" points="281" reactiontime="+122" swimtime="00:08:51.62" resultid="3812" heatid="6485" lane="4" entrytime="00:08:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.36" />
                    <SPLIT distance="100" swimtime="00:02:09.79" />
                    <SPLIT distance="150" swimtime="00:03:22.32" />
                    <SPLIT distance="200" swimtime="00:04:33.37" />
                    <SPLIT distance="250" swimtime="00:05:45.40" />
                    <SPLIT distance="300" swimtime="00:06:57.70" />
                    <SPLIT distance="350" swimtime="00:08:01.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="376" reactiontime="+104" swimtime="00:01:39.63" resultid="3813" heatid="6084" lane="4" entrytime="00:01:44.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="398" reactiontime="+102" swimtime="00:00:45.46" resultid="3814" heatid="6129" lane="5" entrytime="00:00:46.00" entrycourse="SCM" />
                <RESULT eventid="1363" points="256" reactiontime="+90" swimtime="00:00:47.78" resultid="3815" heatid="6225" lane="1" entrytime="00:00:50.00" entrycourse="SCM" />
                <RESULT eventid="1467" points="357" reactiontime="+107" swimtime="00:03:47.10" resultid="3816" heatid="6300" lane="3" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.11" />
                    <SPLIT distance="100" swimtime="00:01:54.45" />
                    <SPLIT distance="150" swimtime="00:03:01.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="287" reactiontime="+120" swimtime="00:04:05.26" resultid="3817" heatid="6373" lane="3" entrytime="00:03:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.20" />
                    <SPLIT distance="100" swimtime="00:02:02.52" />
                    <SPLIT distance="150" swimtime="00:03:09.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="443" reactiontime="+104" swimtime="00:01:43.58" resultid="3818" heatid="6396" lane="3" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-20" firstname="PIOTR" gender="M" lastname="SUWARA" nation="POL" athleteid="3819">
              <RESULTS>
                <RESULT eventid="1137" points="510" swimtime="00:10:23.85" resultid="3820" heatid="6455" lane="6" entrytime="00:10:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.68" />
                    <SPLIT distance="200" swimtime="00:02:30.35" />
                    <SPLIT distance="300" swimtime="00:03:50.22" />
                    <SPLIT distance="400" swimtime="00:05:10.22" />
                    <SPLIT distance="500" swimtime="00:06:29.57" />
                    <SPLIT distance="600" swimtime="00:07:49.91" />
                    <SPLIT distance="700" swimtime="00:09:08.40" />
                    <SPLIT distance="750" swimtime="00:00:03.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="592" reactiontime="+89" swimtime="00:01:00.30" resultid="3821" heatid="6174" lane="3" entrytime="00:01:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="549" reactiontime="+88" swimtime="00:02:16.30" resultid="3822" heatid="6288" lane="3" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:06.28" />
                    <SPLIT distance="150" swimtime="00:01:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="610" reactiontime="+85" swimtime="00:00:27.19" resultid="3823" heatid="6358" lane="1" entrytime="00:00:27.80" entrycourse="SCM" />
                <RESULT eventid="1640" points="527" reactiontime="+92" swimtime="00:04:57.78" resultid="3824" heatid="6567" lane="5" entrytime="00:04:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                    <SPLIT distance="150" swimtime="00:01:46.55" />
                    <SPLIT distance="200" swimtime="00:02:25.16" />
                    <SPLIT distance="250" swimtime="00:03:04.02" />
                    <SPLIT distance="300" swimtime="00:03:42.73" />
                    <SPLIT distance="350" swimtime="00:04:20.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-06-03" firstname="LESZEK" gender="M" lastname="WILKOWSKI" nation="POL" athleteid="3825">
              <RESULTS>
                <RESULT eventid="1137" points="404" swimtime="00:11:39.74" resultid="3826" heatid="6453" lane="6" entrytime="00:11:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.56" />
                    <SPLIT distance="200" swimtime="00:02:46.26" />
                    <SPLIT distance="300" swimtime="00:04:14.28" />
                    <SPLIT distance="400" swimtime="00:05:43.65" />
                    <SPLIT distance="500" swimtime="00:07:14.18" />
                    <SPLIT distance="600" swimtime="00:08:45.58" />
                    <SPLIT distance="700" swimtime="00:10:16.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="394" reactiontime="+92" swimtime="00:00:38.22" resultid="3827" heatid="6132" lane="2" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1302" points="262" reactiontime="+102" swimtime="00:03:23.74" resultid="3828" heatid="6185" lane="3" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                    <SPLIT distance="100" swimtime="00:01:34.94" />
                    <SPLIT distance="150" swimtime="00:02:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="378" reactiontime="+106" swimtime="00:01:23.95" resultid="3829" heatid="6255" lane="2" entrytime="00:01:22.00" entrycourse="SCM" />
                <RESULT eventid="1467" points="463" reactiontime="+99" swimtime="00:02:56.23" resultid="3830" heatid="6305" lane="5" entrytime="00:02:53.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                    <SPLIT distance="100" swimtime="00:01:26.72" />
                    <SPLIT distance="150" swimtime="00:02:18.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="412" reactiontime="+93" swimtime="00:03:02.10" resultid="3831" heatid="6376" lane="2" entrytime="00:03:03.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.83" />
                    <SPLIT distance="100" swimtime="00:02:18.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="407" reactiontime="+94" swimtime="00:01:30.62" resultid="3832" heatid="6401" lane="2" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Grot Koziegłowy" nation="POL">
          <CONTACT name="Ewa Szała" />
          <ATHLETES>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="3834">
              <RESULTS>
                <RESULT eventid="1058" points="710" reactiontime="+99" swimtime="00:06:32.14" resultid="3835" heatid="6431" lane="1" entrytime="00:06:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                    <SPLIT distance="100" swimtime="00:01:31.23" />
                    <SPLIT distance="150" swimtime="00:02:20.24" />
                    <SPLIT distance="200" swimtime="00:03:08.92" />
                    <SPLIT distance="250" swimtime="00:04:04.55" />
                    <SPLIT distance="300" swimtime="00:05:00.38" />
                    <SPLIT distance="350" swimtime="00:05:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="669" reactiontime="+96" swimtime="00:01:26.43" resultid="3836" heatid="6078" lane="2" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="597" reactiontime="+88" swimtime="00:00:41.08" resultid="3837" heatid="6123" lane="6" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1378" points="661" reactiontime="+98" swimtime="00:01:28.65" resultid="3838" heatid="6247" lane="1" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="656" reactiontime="+87" swimtime="00:03:07.74" resultid="3839" heatid="6296" lane="4" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                    <SPLIT distance="100" swimtime="00:01:29.13" />
                    <SPLIT distance="150" swimtime="00:02:23.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="760" reactiontime="+92" swimtime="00:03:07.50" resultid="3840" heatid="6370" lane="2" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.34" />
                    <SPLIT distance="100" swimtime="00:01:32.00" />
                    <SPLIT distance="150" swimtime="00:02:20.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="586" reactiontime="+93" swimtime="00:06:09.27" resultid="3841" heatid="6557" lane="6" entrytime="00:05:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:26.53" />
                    <SPLIT distance="150" swimtime="00:02:13.08" />
                    <SPLIT distance="200" swimtime="00:03:01.73" />
                    <SPLIT distance="250" swimtime="00:03:48.41" />
                    <SPLIT distance="300" swimtime="00:04:35.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Steef Wrocław" nation="POL">
          <CONTACT name="Stefan Skrzypek" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="3843">
              <RESULTS>
                <RESULT eventid="1137" points="595" swimtime="00:11:54.47" resultid="3844" heatid="6451" lane="4" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:12:44.29" />
                    <SPLIT distance="200" swimtime="00:02:54.75" />
                    <SPLIT distance="300" swimtime="00:04:24.08" />
                    <SPLIT distance="400" swimtime="00:05:52.90" />
                    <SPLIT distance="500" swimtime="00:07:23.85" />
                    <SPLIT distance="600" swimtime="00:08:54.82" />
                    <SPLIT distance="700" swimtime="00:10:25.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="436" reactiontime="+96" swimtime="00:03:37.12" resultid="3845" heatid="6111" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.79" />
                    <SPLIT distance="100" swimtime="00:01:45.81" />
                    <SPLIT distance="150" swimtime="00:02:44.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="464" reactiontime="+99" swimtime="00:03:16.59" resultid="3846" heatid="6186" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.61" />
                    <SPLIT distance="100" swimtime="00:01:33.63" />
                    <SPLIT distance="150" swimtime="00:02:25.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="413" reactiontime="+95" swimtime="00:00:37.69" resultid="3847" heatid="6227" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1437" points="582" reactiontime="+106" swimtime="00:02:37.78" resultid="3848" heatid="6283" lane="3" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="100" swimtime="00:01:17.09" />
                    <SPLIT distance="150" swimtime="00:01:57.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="416" reactiontime="+100" swimtime="00:01:26.21" resultid="3849" heatid="6319" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="586" reactiontime="+101" swimtime="00:05:42.01" resultid="3850" heatid="6564" lane="5" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:22.58" />
                    <SPLIT distance="150" swimtime="00:02:06.43" />
                    <SPLIT distance="200" swimtime="00:02:50.73" />
                    <SPLIT distance="250" swimtime="00:03:33.66" />
                    <SPLIT distance="300" swimtime="00:04:16.65" />
                    <SPLIT distance="350" swimtime="00:04:59.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WWSF" name="WOPR Wraszawa SPORT-Figielski" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" email="grzegorz.figielski@sport-figielski.pl" internet="www.sport-figielski.pl" name="Grzegorz Figielski" phone="501294477" state="MAZ" street="Sarmacka 21 m. 41" zip="02-972" />
          <ATHLETES>
            <ATHLETE birthdate="1969-03-04" firstname="Wiktor" gender="M" lastname="Dębski" nation="POL" athleteid="3868">
              <RESULTS>
                <RESULT eventid="1333" points="711" reactiontime="+93" swimtime="00:00:33.04" resultid="3869" heatid="6210" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1363" points="725" reactiontime="+92" swimtime="00:00:29.67" resultid="3870" heatid="6232" lane="6" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Dąbrowa Gornicza" nation="POL" region="SLA">
          <CONTACT name="Waliczek Mariusz" phone="606448210" />
          <ATHLETES>
            <ATHLETE birthdate="1988-03-24" firstname="Kamil" gender="M" lastname="Samul" nation="POL" athleteid="3872">
              <RESULTS>
                <RESULT eventid="1137" points="717" swimtime="00:09:14.10" resultid="3873" heatid="6457" lane="1" entrytime="00:09:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:06.11" />
                    <SPLIT distance="200" swimtime="00:02:15.28" />
                    <SPLIT distance="300" swimtime="00:03:25.16" />
                    <SPLIT distance="400" swimtime="00:04:35.64" />
                    <SPLIT distance="500" swimtime="00:05:45.96" />
                    <SPLIT distance="600" swimtime="00:06:56.96" />
                    <SPLIT distance="700" swimtime="00:08:06.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="843" reactiontime="+80" swimtime="00:01:02.64" resultid="3874" heatid="6099" lane="3" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="718" reactiontime="+76" swimtime="00:00:55.14" resultid="3875" heatid="6180" lane="5" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="713" reactiontime="+79" swimtime="00:02:00.51" resultid="3876" heatid="6292" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:01:00.76" />
                    <SPLIT distance="150" swimtime="00:01:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="685" reactiontime="+75" swimtime="00:00:25.32" resultid="3877" heatid="6365" lane="5" entrytime="00:00:25.00" />
                <RESULT eventid="1640" points="712" reactiontime="+84" swimtime="00:04:20.87" resultid="3878" heatid="6560" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:04.25" />
                    <SPLIT distance="150" swimtime="00:01:37.76" />
                    <SPLIT distance="200" swimtime="00:02:11.19" />
                    <SPLIT distance="250" swimtime="00:02:44.37" />
                    <SPLIT distance="300" swimtime="00:03:17.17" />
                    <SPLIT distance="350" swimtime="00:03:49.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Paweł" gender="M" lastname="Bucki" nation="POL" athleteid="3879">
              <RESULTS>
                <RESULT eventid="1528" points="738" reactiontime="+74" swimtime="00:00:25.16" resultid="3880" heatid="6364" lane="4" entrytime="00:00:25.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Sylwester" gender="M" lastname="Kuster" nation="POL" athleteid="3881">
              <RESULTS>
                <RESULT eventid="1137" points="710" swimtime="00:09:24.84" resultid="3882" heatid="6456" lane="3" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:01:06.35" />
                    <SPLIT distance="200" swimtime="00:02:17.32" />
                    <SPLIT distance="300" swimtime="00:03:28.31" />
                    <SPLIT distance="400" swimtime="00:04:40.35" />
                    <SPLIT distance="500" swimtime="00:05:51.44" />
                    <SPLIT distance="600" swimtime="00:07:03.10" />
                    <SPLIT distance="700" swimtime="00:08:15.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Triathlon Juvenia Wrocław" nation="POL">
          <CONTACT email="maciej.chmura86@gmail.com" name="Chmura" />
          <ATHLETES>
            <ATHLETE birthdate="1986-01-22" firstname="Maciej" gender="M" lastname="Chmura" nation="POL" athleteid="3902">
              <RESULTS>
                <RESULT eventid="1137" points="648" swimtime="00:09:42.23" resultid="6498" heatid="6446" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:10.44" />
                    <SPLIT distance="200" swimtime="00:02:23.40" />
                    <SPLIT distance="300" swimtime="00:03:36.45" />
                    <SPLIT distance="400" swimtime="00:04:49.41" />
                    <SPLIT distance="500" swimtime="00:06:02.25" />
                    <SPLIT distance="600" swimtime="00:07:15.55" />
                    <SPLIT distance="700" swimtime="00:08:28.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="574" reactiontime="+70" swimtime="00:02:13.15" resultid="3904" heatid="6289" lane="2" entrytime="00:02:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:05.79" />
                    <SPLIT distance="150" swimtime="00:01:39.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="3905" heatid="6308" lane="4" entrytime="00:02:40.00" entrycourse="SCM" />
                <RESULT eventid="1640" points="625" reactiontime="+78" swimtime="00:04:42.39" resultid="3906" heatid="6569" lane="1" entrytime="00:04:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:07.43" />
                    <SPLIT distance="150" swimtime="00:01:42.76" />
                    <SPLIT distance="200" swimtime="00:02:18.65" />
                    <SPLIT distance="250" swimtime="00:02:54.39" />
                    <SPLIT distance="300" swimtime="00:03:30.44" />
                    <SPLIT distance="350" swimtime="00:04:06.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MABOL" name="Klub Pływacki Masters Bolesławiec" nation="POL" region="DOL" shortname="Klub Pływacki Masters Bolesław">
          <CONTACT email="sekretarz-masters@o2.pl" name="Marta Satoła" phone="880944737" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="3908">
              <RESULTS>
                <RESULT eventid="1092" points="302" reactiontime="+88" swimtime="00:08:38.68" resultid="3909" heatid="6486" lane="4" entrytime="00:08:22.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.31" />
                    <SPLIT distance="100" swimtime="00:02:04.59" />
                    <SPLIT distance="150" swimtime="00:03:08.47" />
                    <SPLIT distance="200" swimtime="00:04:11.53" />
                    <SPLIT distance="250" swimtime="00:05:25.88" />
                    <SPLIT distance="300" swimtime="00:06:40.72" />
                    <SPLIT distance="350" swimtime="00:07:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="264" reactiontime="+91" swimtime="00:01:52.09" resultid="3910" heatid="6084" lane="2" entrytime="00:01:48.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="181" reactiontime="+93" swimtime="00:04:46.18" resultid="3911" heatid="6185" lane="6" entrytime="00:04:18.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.86" />
                    <SPLIT distance="100" swimtime="00:02:13.39" />
                    <SPLIT distance="150" swimtime="00:03:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="314" reactiontime="+80" swimtime="00:01:48.19" resultid="3912" heatid="6252" lane="1" entrytime="00:01:49.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="269" reactiontime="+90" swimtime="00:04:09.47" resultid="3913" heatid="6300" lane="4" entrytime="00:03:53.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.65" />
                    <SPLIT distance="100" swimtime="00:01:59.01" />
                    <SPLIT distance="150" swimtime="00:03:13.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="164" reactiontime="+85" swimtime="00:02:07.97" resultid="3914" heatid="6317" lane="1" entrytime="00:01:57.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="323" reactiontime="+77" swimtime="00:03:55.92" resultid="3915" heatid="6374" lane="6" entrytime="00:03:48.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.84" />
                    <SPLIT distance="100" swimtime="00:01:55.53" />
                    <SPLIT distance="150" swimtime="00:02:57.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-18" firstname="Marcin" gender="M" lastname="Klimkowski" nation="POL" athleteid="3916">
              <RESULTS>
                <RESULT eventid="1228" points="23" swimtime="00:01:31.61" resultid="3917" heatid="6126" lane="4" entrytime="00:01:39.40" />
                <RESULT eventid="1272" points="11" swimtime="00:03:44.82" resultid="3918" heatid="6159" lane="2" entrytime="00:03:07.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="17" swimtime="00:01:53.24" resultid="3919" heatid="6202" lane="1" entrytime="00:01:52.10" />
                <RESULT eventid="1393" points="26" swimtime="00:03:10.32" resultid="3920" heatid="6250" lane="5" entrytime="00:03:32.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="8" swimtime="00:01:55.04" resultid="3921" heatid="6342" lane="6" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" name="TS Olimpia Poznań" nation="POL" region="WIE">
          <CONTACT name="Pietraszewski Zbigniew" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="3929">
              <RESULTS>
                <RESULT eventid="1257" points="515" reactiontime="+96" swimtime="00:01:29.05" resultid="3930" heatid="6151" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="437" reactiontime="+101" swimtime="00:00:50.84" resultid="3931" heatid="6196" lane="6" entrytime="00:00:52.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="3932" heatid="6274" lane="5" entrytime="00:03:20.00" />
                <RESULT eventid="1513" points="614" reactiontime="+100" swimtime="00:00:37.81" resultid="3933" heatid="6333" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1595" points="452" reactiontime="+104" swimtime="00:01:52.62" resultid="3934" heatid="6506" lane="1" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Grażyna" gender="F" lastname="Cabaj-Drela" nation="POL" athleteid="3935">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. G" eventid="1183" points="871" reactiontime="+92" swimtime="00:03:18.81" resultid="3936" heatid="6105" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                    <SPLIT distance="100" swimtime="00:01:34.53" />
                    <SPLIT distance="150" swimtime="00:02:26.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="734" reactiontime="+91" swimtime="00:00:42.64" resultid="3937" heatid="6198" lane="1" entrytime="00:00:45.00" />
                <RESULT comment="Rekord Polski kat. G" eventid="1378" points="829" reactiontime="+80" swimtime="00:01:27.25" resultid="3938" heatid="6246" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="808" reactiontime="+90" swimtime="00:01:33.73" resultid="3939" heatid="6508" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="Lesiński" nation="POL" athleteid="3940">
              <RESULTS>
                <RESULT eventid="1168" points="521" reactiontime="+114" swimtime="00:01:33.89" resultid="3941" heatid="6086" lane="1" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="577" reactiontime="+79" swimtime="00:00:42.36" resultid="3942" heatid="6130" lane="1" entrytime="00:00:44.00" />
                <RESULT eventid="1393" points="538" reactiontime="+77" swimtime="00:01:38.30" resultid="3943" heatid="6253" lane="1" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="3944" heatid="6301" lane="3" entrytime="00:03:38.00" />
                <RESULT eventid="1558" points="497" reactiontime="+81" swimtime="00:03:40.31" resultid="3945" heatid="6374" lane="4" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.58" />
                    <SPLIT distance="100" swimtime="00:01:44.74" />
                    <SPLIT distance="150" swimtime="00:02:42.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Janusz" gender="M" lastname="Woch" nation="POL" athleteid="3946">
              <RESULTS>
                <RESULT eventid="1092" points="483" reactiontime="+87" swimtime="00:07:56.43" resultid="3947" heatid="6486" lane="3" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.86" />
                    <SPLIT distance="100" swimtime="00:02:01.18" />
                    <SPLIT distance="150" swimtime="00:03:01.95" />
                    <SPLIT distance="200" swimtime="00:04:00.17" />
                    <SPLIT distance="250" swimtime="00:05:00.03" />
                    <SPLIT distance="300" swimtime="00:05:59.98" />
                    <SPLIT distance="350" swimtime="00:06:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="531" reactiontime="+91" swimtime="00:01:33.27" resultid="3948" heatid="6086" lane="2" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="575" reactiontime="+79" swimtime="00:03:41.91" resultid="3949" heatid="6111" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.31" />
                    <SPLIT distance="100" swimtime="00:01:47.52" />
                    <SPLIT distance="150" swimtime="00:02:46.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="588" reactiontime="+82" swimtime="00:00:43.19" resultid="3950" heatid="6208" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1393" points="491" reactiontime="+83" swimtime="00:01:41.32" resultid="3951" heatid="6253" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="564" reactiontime="+96" swimtime="00:03:31.20" resultid="3952" heatid="6375" lane="1" entrytime="00:03:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.15" />
                    <SPLIT distance="100" swimtime="00:01:40.75" />
                    <SPLIT distance="150" swimtime="00:02:36.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="553" reactiontime="+85" swimtime="00:01:39.17" resultid="3953" heatid="6398" lane="4" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="3954">
              <RESULTS>
                <RESULT eventid="1137" points="323" swimtime="00:14:44.72" resultid="3955" heatid="6449" lane="6" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.39" />
                    <SPLIT distance="200" swimtime="00:03:31.04" />
                    <SPLIT distance="300" swimtime="00:05:22.41" />
                    <SPLIT distance="400" swimtime="00:07:12.38" />
                    <SPLIT distance="500" swimtime="00:09:05.70" />
                    <SPLIT distance="600" swimtime="00:11:01.57" />
                    <SPLIT distance="700" swimtime="00:12:55.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="556" reactiontime="+76" swimtime="00:00:40.66" resultid="3956" heatid="6130" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1393" points="465" reactiontime="+74" swimtime="00:01:34.98" resultid="3957" heatid="6253" lane="4" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="3958" heatid="6375" lane="6" entrytime="00:03:32.00" />
                <RESULT eventid="1640" points="353" reactiontime="+104" swimtime="00:06:57.47" resultid="3959" heatid="6561" lane="3" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                    <SPLIT distance="100" swimtime="00:01:39.15" />
                    <SPLIT distance="150" swimtime="00:02:32.50" />
                    <SPLIT distance="200" swimtime="00:03:26.02" />
                    <SPLIT distance="250" swimtime="00:04:20.33" />
                    <SPLIT distance="300" swimtime="00:05:14.20" />
                    <SPLIT distance="350" swimtime="00:06:07.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="3960">
              <RESULTS>
                <RESULT eventid="1092" points="597" reactiontime="+90" swimtime="00:06:41.30" resultid="3961" heatid="6488" lane="3" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.17" />
                    <SPLIT distance="100" swimtime="00:01:41.99" />
                    <SPLIT distance="150" swimtime="00:02:30.46" />
                    <SPLIT distance="200" swimtime="00:03:18.90" />
                    <SPLIT distance="250" swimtime="00:04:14.92" />
                    <SPLIT distance="300" swimtime="00:05:09.05" />
                    <SPLIT distance="350" swimtime="00:05:56.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="531" reactiontime="+90" swimtime="00:01:23.96" resultid="3962" heatid="6090" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="459" reactiontime="+82" swimtime="00:00:41.35" resultid="3963" heatid="6132" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1393" points="460" reactiontime="+74" swimtime="00:01:27.48" resultid="3964" heatid="6255" lane="6" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="590" reactiontime="+90" swimtime="00:03:04.51" resultid="3965" heatid="6304" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:30.53" />
                    <SPLIT distance="150" swimtime="00:02:22.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="544" reactiontime="+80" swimtime="00:03:04.42" resultid="3966" heatid="6376" lane="3" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:01:30.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="3967">
              <RESULTS>
                <RESULT eventid="1198" points="691" reactiontime="+79" swimtime="00:02:54.16" resultid="3968" heatid="6115" lane="5" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                    <SPLIT distance="100" swimtime="00:01:25.17" />
                    <SPLIT distance="150" swimtime="00:02:10.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="645" reactiontime="+81" swimtime="00:01:03.39" resultid="3969" heatid="6171" lane="5" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="631" reactiontime="+81" swimtime="00:00:35.80" resultid="3970" heatid="6214" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="3971" heatid="6287" lane="1" entrytime="00:02:23.00" />
                <RESULT eventid="1610" points="684" reactiontime="+78" swimtime="00:01:18.00" resultid="3972" heatid="6406" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Radosław" gender="M" lastname="Pierz" nation="POL" athleteid="3973">
              <RESULTS>
                <RESULT eventid="1168" points="320" reactiontime="+91" swimtime="00:01:30.17" resultid="3974" heatid="6087" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="366" reactiontime="+85" swimtime="00:00:41.23" resultid="3975" heatid="6208" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1363" points="231" reactiontime="+99" swimtime="00:00:43.45" resultid="3976" heatid="6226" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1528" points="366" reactiontime="+91" swimtime="00:00:34.12" resultid="3977" heatid="6346" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1610" points="340" reactiontime="+90" swimtime="00:01:36.21" resultid="3978" heatid="6399" lane="6" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Łukasz" gender="M" lastname="Bogucki" nation="POL" athleteid="3979">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="3980" heatid="6094" lane="6" entrytime="00:01:13.00" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="3981" heatid="6136" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1363" status="DNS" swimtime="00:00:00.00" resultid="3982" heatid="6236" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="3983" heatid="6356" lane="4" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+80" swimtime="00:02:45.48" resultid="3985" heatid="6524" lane="1" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                    <SPLIT distance="100" swimtime="00:01:25.24" />
                    <SPLIT distance="150" swimtime="00:02:07.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3954" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3946" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="3960" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3940" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+85" swimtime="00:02:15.23" resultid="3986" heatid="6496" lane="1" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                    <SPLIT distance="100" swimtime="00:01:03.58" />
                    <SPLIT distance="150" swimtime="00:01:36.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3967" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="3935" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3960" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3929" number="4" reactiontime="+81" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ORSOPOLE" name="Odrzańskie Ratownictwo Specjalistyczne Opole" nation="POL" region="OPO" shortname="Odrzańskie Ratownictwo Specjal">
          <CONTACT email="wkania62@gmail.com" name="Kania" />
          <ATHLETES>
            <ATHLETE birthdate="1973-01-01" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="3994">
              <RESULTS>
                <RESULT eventid="1153" points="494" reactiontime="+98" swimtime="00:01:25.61" resultid="3995" heatid="6079" lane="5" entrytime="00:01:26.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="474" reactiontime="+72" swimtime="00:00:40.15" resultid="3996" heatid="6123" lane="2" entrytime="00:00:40.25" />
                <RESULT eventid="1378" points="410" reactiontime="+77" swimtime="00:01:27.10" resultid="3997" heatid="6247" lane="6" entrytime="00:01:26.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="414" reactiontime="+108" swimtime="00:03:10.61" resultid="3998" heatid="6295" lane="3" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:29.84" />
                    <SPLIT distance="150" swimtime="00:02:25.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="399" reactiontime="+72" swimtime="00:03:07.98" resultid="3999" heatid="6369" lane="3" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                    <SPLIT distance="100" swimtime="00:01:30.30" />
                    <SPLIT distance="150" swimtime="00:02:20.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Grzegorz" gender="M" lastname="Stanek" nation="POL" athleteid="4000">
              <RESULTS>
                <RESULT eventid="1092" points="869" reactiontime="+85" swimtime="00:05:07.39" resultid="4001" heatid="6492" lane="4" entrytime="00:05:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                    <SPLIT distance="150" swimtime="00:01:49.44" />
                    <SPLIT distance="200" swimtime="00:02:28.34" />
                    <SPLIT distance="250" swimtime="00:03:12.57" />
                    <SPLIT distance="300" swimtime="00:03:56.88" />
                    <SPLIT distance="350" swimtime="00:04:32.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Wojciech" gender="M" lastname="Stanek" nation="POL" athleteid="4002">
              <RESULTS>
                <RESULT eventid="1092" points="433" reactiontime="+70" swimtime="00:05:49.07" resultid="4003" heatid="6491" lane="1" entrytime="00:05:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:01:24.87" />
                    <SPLIT distance="150" swimtime="00:02:10.14" />
                    <SPLIT distance="200" swimtime="00:02:54.61" />
                    <SPLIT distance="250" swimtime="00:03:41.08" />
                    <SPLIT distance="300" swimtime="00:04:28.29" />
                    <SPLIT distance="350" swimtime="00:05:09.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Waldemar" gender="M" lastname="Kania" nation="POL" athleteid="4004">
              <RESULTS>
                <RESULT eventid="1437" points="526" reactiontime="+92" swimtime="00:02:33.92" resultid="4007" heatid="6285" lane="1" entrytime="00:02:32.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:14.02" />
                    <SPLIT distance="150" swimtime="00:01:54.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="4008" heatid="6379" lane="2" entrytime="00:02:40.11" />
                <RESULT eventid="1137" points="584" swimtime="00:11:18.22" resultid="4005" heatid="6453" lane="2" entrytime="00:11:20.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:20.19" />
                    <SPLIT distance="200" swimtime="00:02:45.18" />
                    <SPLIT distance="300" swimtime="00:04:10.22" />
                    <SPLIT distance="400" swimtime="00:05:35.32" />
                    <SPLIT distance="500" swimtime="00:07:01.33" />
                    <SPLIT distance="600" swimtime="00:08:27.62" />
                    <SPLIT distance="700" swimtime="00:09:53.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="542" reactiontime="+97" swimtime="00:01:09.75" resultid="4006" heatid="6168" lane="1" entrytime="00:01:09.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="537" reactiontime="+97" swimtime="00:05:30.02" resultid="6572" heatid="6567" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                    <SPLIT distance="100" swimtime="00:01:18.55" />
                    <SPLIT distance="150" swimtime="00:02:00.60" />
                    <SPLIT distance="200" swimtime="00:02:42.88" />
                    <SPLIT distance="250" swimtime="00:03:24.93" />
                    <SPLIT distance="300" swimtime="00:04:07.38" />
                    <SPLIT distance="350" swimtime="00:04:49.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Marcin" gender="M" lastname="Wilczyński" nation="POL" athleteid="4010">
              <RESULTS>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="4011" heatid="6115" lane="3" entrytime="00:02:50.65" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="4012" heatid="6214" lane="5" entrytime="00:00:34.65" />
                <RESULT eventid="1610" points="776" reactiontime="+89" swimtime="00:01:13.09" resultid="4013" heatid="6406" lane="2" entrytime="00:01:17.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Grzegorz" gender="M" lastname="Bielaczyc" nation="POL" athleteid="4014">
              <RESULTS>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="4015" heatid="6210" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1363" status="DNS" swimtime="00:00:00.00" resultid="4016" heatid="6226" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Stowarzyszenie Pływackie &quot;Swimmers&quot;Warszawa" nation="POL" region="MAZ" shortname="Stowarzyszenie Pływackie &quot;Swim">
          <CONTACT city="WARSZAWA" email="info@swimmersteam.pl" internet="www.swimmersteam.pl" name="REMIGIUSZ GOŁĘBIOWSKI" phone="601333782" state="MAZ" street="GŁADKA 18" zip="02-172" />
          <ATHLETES>
            <ATHLETE birthdate="1984-12-07" firstname="Margarita" gender="F" lastname="Aragon de Szumańska" nation="POL" athleteid="4018">
              <RESULTS>
                <RESULT eventid="1213" points="335" reactiontime="+83" swimtime="00:00:43.83" resultid="4019" heatid="6123" lane="3" entrytime="00:00:39.00" entrycourse="SCM" />
                <RESULT eventid="1513" points="413" reactiontime="+83" swimtime="00:00:35.44" resultid="4020" heatid="6336" lane="6" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1625" reactiontime="+117" status="DNS" swimtime="00:00:00.00" resultid="4021" heatid="6556" lane="3" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:01:29.20" />
                    <SPLIT distance="150" swimtime="00:02:19.29" />
                    <SPLIT distance="200" swimtime="00:03:10.78" />
                    <SPLIT distance="250" swimtime="00:04:00.78" />
                    <SPLIT distance="300" swimtime="00:04:53.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-07-07" firstname="REMIGIUSZ" gender="M" lastname="GOŁĘBIOWSKI" nation="POL" athleteid="4022">
              <RESULTS>
                <RESULT eventid="1168" points="646" reactiontime="+77" swimtime="00:01:07.54" resultid="4023" heatid="6097" lane="2" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="632" reactiontime="+73" swimtime="00:00:59.90" resultid="4024" heatid="6178" lane="6" entrytime="00:00:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="4025" heatid="6214" lane="3" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1363" points="679" reactiontime="+80" swimtime="00:00:28.59" resultid="4026" heatid="6241" lane="6" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="1498" points="639" reactiontime="+79" swimtime="00:01:06.24" resultid="4027" heatid="6326" lane="6" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="640" reactiontime="+81" swimtime="00:00:26.86" resultid="4028" heatid="6360" lane="2" entrytime="00:00:26.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="Redeco Wrocław" nation="POL" region="DOL">
          <CONTACT city="Wrocław" name="Wolny Dariusz" phone="603630870" state="DOL" street="Rogowska 52a" zip="54-440" />
          <ATHLETES>
            <ATHLETE birthdate="1960-03-21" firstname="Dariusz" gender="M" lastname="Wolny" nation="POL" athleteid="4030">
              <RESULTS>
                <RESULT eventid="1168" points="966" reactiontime="+77" swimtime="00:01:06.27" resultid="4031" heatid="6097" lane="1" entrytime="00:01:07.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="1014" reactiontime="+61" swimtime="00:00:30.47" resultid="4032" heatid="6137" lane="5" entrytime="00:00:30.77" />
                <RESULT eventid="1393" points="1024" reactiontime="+70" swimtime="00:01:06.64" resultid="4033" heatid="6261" lane="1" entrytime="00:01:07.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="4034" heatid="6310" lane="4" entrytime="00:02:25.77" />
                <RESULT eventid="1558" points="1092" reactiontime="+70" swimtime="00:02:24.65" resultid="4035" heatid="6381" lane="3" entrytime="00:02:25.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:10.19" />
                    <SPLIT distance="150" swimtime="00:01:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="843" reactiontime="+79" swimtime="00:01:17.03" resultid="4036" heatid="6406" lane="5" entrytime="00:01:17.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Joanna" gender="F" lastname="Chojcan" nation="POL" athleteid="4037">
              <RESULTS>
                <RESULT eventid="1058" points="575" reactiontime="+77" swimtime="00:06:04.27" resultid="4038" heatid="6431" lane="4" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:19.18" />
                    <SPLIT distance="150" swimtime="00:02:05.36" />
                    <SPLIT distance="200" swimtime="00:02:51.26" />
                    <SPLIT distance="250" swimtime="00:03:44.20" />
                    <SPLIT distance="300" swimtime="00:04:37.79" />
                    <SPLIT distance="350" swimtime="00:05:21.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="625" reactiontime="+65" swimtime="00:00:35.61" resultid="4039" heatid="6125" lane="1" entrytime="00:00:35.90" />
                <RESULT eventid="1287" points="444" reactiontime="+83" swimtime="00:03:02.07" resultid="4040" heatid="6182" lane="4" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:01:23.46" />
                    <SPLIT distance="150" swimtime="00:02:11.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="533" reactiontime="+65" swimtime="00:01:18.25" resultid="4041" heatid="6248" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="564" reactiontime="+81" swimtime="00:02:51.82" resultid="4042" heatid="6297" lane="4" entrytime="00:02:53.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:18.36" />
                    <SPLIT distance="150" swimtime="00:02:10.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="494" reactiontime="+80" swimtime="00:01:19.88" resultid="4043" heatid="6315" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="494" reactiontime="+70" swimtime="00:02:50.96" resultid="4044" heatid="6371" lane="1" entrytime="00:02:51.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:01:21.55" />
                    <SPLIT distance="150" swimtime="00:02:06.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-25" firstname="Marlena" gender="F" lastname="Jakubów" nation="POL" athleteid="4045">
              <RESULTS>
                <RESULT eventid="1058" points="314" reactiontime="+106" swimtime="00:07:36.99" resultid="4046" heatid="6430" lane="2" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.62" />
                    <SPLIT distance="100" swimtime="00:01:49.94" />
                    <SPLIT distance="150" swimtime="00:02:50.26" />
                    <SPLIT distance="200" swimtime="00:03:53.02" />
                    <SPLIT distance="250" swimtime="00:04:53.19" />
                    <SPLIT distance="300" swimtime="00:05:55.22" />
                    <SPLIT distance="350" swimtime="00:06:47.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="345" reactiontime="+94" swimtime="00:00:44.60" resultid="4047" heatid="6121" lane="4" entrytime="00:00:45.87" />
                <RESULT eventid="1257" points="357" reactiontime="+114" swimtime="00:01:21.35" resultid="4048" heatid="6152" lane="2" entrytime="00:01:25.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="213" reactiontime="+97" swimtime="00:01:48.34" resultid="4049" heatid="6245" lane="1" entrytime="00:01:47.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="288" reactiontime="+105" swimtime="00:03:10.42" resultid="4050" heatid="6274" lane="3" entrytime="00:03:09.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.75" />
                    <SPLIT distance="100" swimtime="00:02:23.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="424" reactiontime="+106" swimtime="00:00:35.65" resultid="4051" heatid="6335" lane="5" entrytime="00:00:35.72" />
                <RESULT eventid="1543" points="225" reactiontime="+100" swimtime="00:03:47.39" resultid="4052" heatid="6368" lane="1" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.78" />
                    <SPLIT distance="100" swimtime="00:01:50.81" />
                    <SPLIT distance="150" swimtime="00:02:51.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-27" firstname="Hanna" gender="F" lastname="Sikacz" nation="POL" athleteid="4053">
              <RESULTS>
                <RESULT eventid="1122" points="452" swimtime="00:12:16.58" resultid="4054" heatid="6444" lane="2" entrytime="00:12:03.97">
                  <SPLITS>
                    <SPLIT distance="400" swimtime="00:06:04.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="374" reactiontime="+86" swimtime="00:01:30.19" resultid="4055" heatid="6079" lane="1" entrytime="00:01:27.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="420" reactiontime="+83" swimtime="00:01:17.51" resultid="4056" heatid="6154" lane="1" entrytime="00:01:17.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="411" reactiontime="+88" swimtime="00:02:48.40" resultid="4057" heatid="6276" lane="1" entrytime="00:02:48.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:20.01" />
                    <SPLIT distance="150" swimtime="00:02:05.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="393" reactiontime="+80" swimtime="00:03:15.06" resultid="4058" heatid="6296" lane="6" entrytime="00:03:12.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.60" />
                    <SPLIT distance="100" swimtime="00:01:37.08" />
                    <SPLIT distance="150" swimtime="00:02:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="280" reactiontime="+80" swimtime="00:01:37.75" resultid="4059" heatid="6314" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="432" reactiontime="+80" swimtime="00:05:54.64" resultid="4060" heatid="6557" lane="1" entrytime="00:05:46.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:02:08.21" />
                    <SPLIT distance="200" swimtime="00:02:53.18" />
                    <SPLIT distance="250" swimtime="00:03:39.23" />
                    <SPLIT distance="300" swimtime="00:04:25.44" />
                    <SPLIT distance="350" swimtime="00:05:11.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-23" firstname="Agnieszka" gender="F" lastname="Bystrzycka" nation="POL" athleteid="4061">
              <RESULTS>
                <RESULT eventid="1183" points="862" reactiontime="+82" swimtime="00:02:42.99" resultid="4062" heatid="6107" lane="3" entrytime="00:02:39.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:16.77" />
                    <SPLIT distance="150" swimtime="00:01:59.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="952" reactiontime="+78" swimtime="00:00:33.83" resultid="4063" heatid="6201" lane="3" entrytime="00:00:33.97" />
                <RESULT eventid="1595" points="878" reactiontime="+80" swimtime="00:01:14.54" resultid="4064" heatid="6510" lane="3" entrytime="00:01:14.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Dariusz" gender="M" lastname="Patrzałek" nation="POL" athleteid="4065">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="4066" heatid="6084" lane="5" entrytime="00:01:48.85" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="4068" heatid="6204" lane="6" entrytime="00:00:52.52" />
                <RESULT eventid="1363" status="DNS" swimtime="00:00:00.00" resultid="4069" heatid="6226" lane="6" entrytime="00:00:44.63" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="4070" heatid="6343" lane="3" entrytime="00:00:39.90" />
                <RESULT eventid="1610" status="DNS" swimtime="00:00:00.00" resultid="4071" heatid="6396" lane="2" entrytime="00:01:50.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-28" firstname="Przemysław" gender="M" lastname="Matuszek" nation="POL" athleteid="4072">
              <RESULTS>
                <RESULT eventid="1168" points="481" reactiontime="+83" swimtime="00:01:14.37" resultid="4073" heatid="6093" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="401" reactiontime="+79" swimtime="00:01:08.63" resultid="4074" heatid="6172" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="550" reactiontime="+80" swimtime="00:00:30.82" resultid="4075" heatid="6236" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="4076" heatid="6287" lane="6" entrytime="00:02:25.00" />
                <RESULT eventid="1498" points="414" reactiontime="+81" swimtime="00:01:14.71" resultid="4077" heatid="6323" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" status="DNS" swimtime="00:00:00.00" resultid="4078" heatid="6403" lane="1" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-07" firstname="Wojciech" gender="M" lastname="Ducki" nation="POL" athleteid="4079">
              <RESULTS>
                <RESULT eventid="1168" points="581" reactiontime="+74" swimtime="00:01:16.19" resultid="4080" heatid="6091" lane="2" entrytime="00:01:18.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="601" reactiontime="+77" swimtime="00:01:04.89" resultid="4081" heatid="6170" lane="1" entrytime="00:01:05.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="599" reactiontime="+65" swimtime="00:00:32.48" resultid="4082" heatid="6232" lane="2" entrytime="00:00:31.91" />
                <RESULT comment="O4 - przedwczesny start." eventid="1528" reactiontime="+43" status="DSQ" swimtime="00:00:28.57" resultid="4083" heatid="6355" lane="5" entrytime="00:00:28.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-03-16" firstname="Katarzyna" gender="F" lastname="Krawczyk" nation="POL" athleteid="4084">
              <RESULTS>
                <RESULT eventid="1153" points="422" reactiontime="+76" swimtime="00:01:27.41" resultid="4085" heatid="6081" lane="4" entrytime="00:01:18.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="408" reactiontime="+78" swimtime="00:01:17.41" resultid="4086" heatid="6155" lane="1" entrytime="00:01:14.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="4087" heatid="6197" lane="3" entrytime="00:00:47.47" />
                <RESULT eventid="1348" points="517" reactiontime="+77" swimtime="00:00:36.30" resultid="4088" heatid="6220" lane="4" entrytime="00:00:38.58" />
                <RESULT eventid="1483" points="311" reactiontime="+80" swimtime="00:01:33.14" resultid="4089" heatid="6314" lane="4" entrytime="00:01:33.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="468" reactiontime="+79" swimtime="00:00:34.00" resultid="4090" heatid="6335" lane="4" entrytime="00:00:35.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-10" firstname="Maciej" gender="M" lastname="Koszarek" nation="POL" athleteid="4091">
              <RESULTS>
                <RESULT eventid="1272" points="447" reactiontime="+104" swimtime="00:01:06.13" resultid="4093" heatid="6166" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="4094" heatid="6186" lane="4" entrytime="00:03:20.00" />
                <RESULT eventid="1363" points="502" reactiontime="+88" swimtime="00:00:31.89" resultid="4095" heatid="6233" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1437" points="379" reactiontime="+96" swimtime="00:02:32.87" resultid="4096" heatid="6286" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:12.71" />
                    <SPLIT distance="150" swimtime="00:01:53.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="404" reactiontime="+97" swimtime="00:01:15.10" resultid="4097" heatid="6320" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="412" reactiontime="+86" swimtime="00:00:30.56" resultid="4098" heatid="6353" lane="6" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-26" firstname="Wojciech" gender="M" lastname="Urban" nation="POL" athleteid="4099">
              <RESULTS>
                <RESULT eventid="1272" points="710" reactiontime="+78" swimtime="00:00:56.76" resultid="4100" heatid="6177" lane="1" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="705" reactiontime="+81" swimtime="00:00:28.38" resultid="4101" heatid="6238" lane="3" entrytime="00:00:28.99" />
                <RESULT eventid="1528" points="770" reactiontime="+77" swimtime="00:00:25.16" resultid="4102" heatid="6364" lane="5" entrytime="00:00:25.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-01" firstname="Wojciech" gender="M" lastname="Dobrowolski" nation="POL" athleteid="4103">
              <RESULTS>
                <RESULT eventid="1168" points="414" reactiontime="+87" swimtime="00:01:17.66" resultid="4104" heatid="6090" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="469" reactiontime="+84" swimtime="00:01:05.06" resultid="4105" heatid="6169" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="452" reactiontime="+90" swimtime="00:00:33.03" resultid="4106" heatid="6230" lane="5" entrytime="00:00:33.33" />
                <RESULT eventid="1437" points="393" reactiontime="+97" swimtime="00:02:31.03" resultid="4107" heatid="6286" lane="5" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:13.10" />
                    <SPLIT distance="150" swimtime="00:01:54.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="490" reactiontime="+86" swimtime="00:00:28.84" resultid="4108" heatid="6355" lane="3" entrytime="00:00:28.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-12-13" firstname="Agata" gender="F" lastname="Grochowska" nation="POL" athleteid="4109">
              <RESULTS>
                <RESULT eventid="1122" points="223" swimtime="00:15:33.33" resultid="4110" heatid="6444" lane="4" entrytime="00:12:00.00" />
                <RESULT comment="Zmiana stylu." eventid="1153" reactiontime="+90" status="DSQ" swimtime="00:01:41.35" resultid="4111" heatid="6077" lane="6" entrytime="00:01:44.00" />
                <RESULT eventid="1213" points="336" reactiontime="+71" swimtime="00:00:45.21" resultid="4112" heatid="6121" lane="1" entrytime="00:00:49.00" />
                <RESULT eventid="1318" points="373" reactiontime="+89" swimtime="00:00:47.23" resultid="4113" heatid="6196" lane="1" entrytime="00:00:51.00" />
                <RESULT eventid="1378" points="310" reactiontime="+63" swimtime="00:01:38.50" resultid="4114" heatid="6245" lane="5" entrytime="00:01:36.55" />
                <RESULT eventid="1513" points="360" reactiontime="+89" swimtime="00:00:38.22" resultid="4115" heatid="6333" lane="3" entrytime="00:00:37.36" />
                <RESULT eventid="1543" points="299" reactiontime="+71" swimtime="00:03:37.48" resultid="4116" heatid="6370" lane="5" entrytime="00:03:08.08">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:40.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+75" swimtime="00:01:48.69" resultid="4120" heatid="6533" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                    <SPLIT distance="100" swimtime="00:00:56.72" />
                    <SPLIT distance="150" swimtime="00:01:23.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4079" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4072" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="4030" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4099" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+62" swimtime="00:02:03.45" resultid="4118" heatid="6524" lane="4" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:06.71" />
                    <SPLIT distance="150" swimtime="00:01:38.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4030" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4072" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="4079" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="4099" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1243" reactiontime="+70" swimtime="00:02:20.20" resultid="4119" heatid="6520" lane="3" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                    <SPLIT distance="100" swimtime="00:01:09.50" />
                    <SPLIT distance="150" swimtime="00:01:45.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4037" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4061" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="4084" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4053" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1408" reactiontime="+80" swimtime="00:02:07.32" resultid="4121" heatid="6528" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                    <SPLIT distance="100" swimtime="00:01:03.08" />
                    <SPLIT distance="150" swimtime="00:01:36.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4061" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4037" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="4084" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4053" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+76" swimtime="00:02:29.97" resultid="4124" heatid="6537" lane="4" entrytime="00:02:15.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:29.53" />
                    <SPLIT distance="150" swimtime="00:02:01.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4091" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4053" number="2" reactiontime="-50" />
                    <RELAYPOSITION athleteid="4045" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4103" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+81" swimtime="00:02:06.97" resultid="4125" heatid="6497" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                    <SPLIT distance="100" swimtime="00:00:58.53" />
                    <SPLIT distance="150" swimtime="00:01:38.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4079" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4030" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="4053" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="4045" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+78" swimtime="00:01:54.06" resultid="4117" heatid="6497" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                    <SPLIT distance="100" swimtime="00:01:00.43" />
                    <SPLIT distance="150" swimtime="00:01:28.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4061" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4103" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="4084" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="4099" number="4" reactiontime="+92" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+68" swimtime="00:02:16.52" resultid="4122" heatid="6538" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4030" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4072" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="4084" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4037" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+82" swimtime="00:02:08.16" resultid="4123" heatid="6497" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.33" />
                    <SPLIT distance="150" swimtime="00:01:38.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4091" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="4072" number="2" />
                    <RELAYPOSITION athleteid="4037" number="3" reactiontime="+1" />
                    <RELAYPOSITION athleteid="4109" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Weteran Zabrze" nation="POL">
          <CONTACT city="ZABRZE" name="BOSOWSKI WŁODZIMIERZ" street="ŚW.JANA  4 A/4" zip="41803" />
          <ATHLETES>
            <ATHLETE birthdate="1986-01-01" firstname="Krzysztof" gender="M" lastname="Nowak" nation="POL" athleteid="3859">
              <RESULTS>
                <RESULT eventid="1272" points="655" reactiontime="+71" swimtime="00:00:58.22" resultid="3860" heatid="6175" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="730" reactiontime="+73" swimtime="00:00:28.16" resultid="3861" heatid="6237" lane="3" entrytime="00:00:29.60" />
                <RESULT eventid="1528" points="667" reactiontime="+70" swimtime="00:00:26.02" resultid="3862" heatid="6363" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="1640" points="534" reactiontime="+72" swimtime="00:04:57.50" resultid="3863" heatid="6568" lane="1" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:08.20" />
                    <SPLIT distance="150" swimtime="00:01:45.16" />
                    <SPLIT distance="200" swimtime="00:02:23.67" />
                    <SPLIT distance="250" swimtime="00:03:02.06" />
                    <SPLIT distance="300" swimtime="00:03:41.17" />
                    <SPLIT distance="350" swimtime="00:04:19.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="GENOWEFA" gender="F" lastname="DRUŻYŃSKA" nation="POL" athleteid="4137">
              <RESULTS>
                <RESULT eventid="1318" points="383" swimtime="00:00:53.13" resultid="4138" heatid="6194" lane="2" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="ALFRED" gender="M" lastname="ZABRZAŃSKI" nation="POL" athleteid="4139">
              <RESULTS>
                <RESULT eventid="1137" points="520" swimtime="00:12:27.14" resultid="4140" heatid="6450" lane="1" entrytime="00:12:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                    <SPLIT distance="100" swimtime="00:01:24.00" />
                    <SPLIT distance="200" swimtime="00:02:54.60" />
                    <SPLIT distance="300" swimtime="00:04:27.41" />
                    <SPLIT distance="400" swimtime="00:06:02.04" />
                    <SPLIT distance="500" swimtime="00:07:38.56" />
                    <SPLIT distance="600" swimtime="00:09:14.81" />
                    <SPLIT distance="700" swimtime="00:10:51.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="544" reactiontime="+83" swimtime="00:01:23.31" resultid="4141" heatid="6087" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="645" reactiontime="+77" swimtime="00:01:07.90" resultid="4142" heatid="6168" lane="6" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="573" reactiontime="+91" swimtime="00:02:38.65" resultid="4143" heatid="6283" lane="6" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:14.57" />
                    <SPLIT distance="150" swimtime="00:01:56.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="605" reactiontime="+73" swimtime="00:00:30.86" resultid="4144" heatid="6351" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="1640" points="539" reactiontime="+90" swimtime="00:05:51.78" resultid="4145" heatid="6563" lane="2" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:23.36" />
                    <SPLIT distance="150" swimtime="00:02:08.85" />
                    <SPLIT distance="200" swimtime="00:02:56.47" />
                    <SPLIT distance="250" swimtime="00:03:43.71" />
                    <SPLIT distance="300" swimtime="00:04:29.59" />
                    <SPLIT distance="350" swimtime="00:05:13.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="AURELIA" gender="F" lastname="WRONA" nation="POL" athleteid="4146">
              <RESULTS>
                <RESULT eventid="1213" points="617" reactiontime="+73" swimtime="00:00:43.51" resultid="4147" heatid="6122" lane="4" entrytime="00:00:43.00" />
                <RESULT eventid="1378" points="651" reactiontime="+79" swimtime="00:01:34.56" resultid="4148" heatid="6246" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="509" reactiontime="+88" swimtime="00:00:38.85" resultid="4149" heatid="6335" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1543" points="711" reactiontime="+78" swimtime="00:03:27.79" resultid="4150" heatid="6369" lane="1" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                    <SPLIT distance="100" swimtime="00:01:42.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="MARIA" gender="F" lastname="BUCZKOWSKA" nation="POL" athleteid="4151">
              <RESULTS>
                <RESULT eventid="1183" points="740" reactiontime="+110" swimtime="00:03:59.19" resultid="4152" heatid="6104" lane="6" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="766" swimtime="00:00:47.90" resultid="4153" heatid="6197" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="1595" points="702" reactiontime="+102" swimtime="00:01:49.39" resultid="4154" heatid="6506" lane="6" entrytime="00:01:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-01-01" firstname="WŁADYSŁAW" gender="M" lastname="BUCZKOWSKI" nation="POL" athleteid="4155">
              <RESULTS>
                <RESULT eventid="1228" points="651" reactiontime="+83" swimtime="00:00:44.08" resultid="4156" heatid="6129" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1272" points="597" reactiontime="+90" swimtime="00:01:19.63" resultid="4157" heatid="6162" lane="3" entrytime="00:01:16.00" />
                <RESULT eventid="1333" points="879" reactiontime="+73" swimtime="00:00:39.90" resultid="4158" heatid="6210" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1437" points="592" reactiontime="+107" swimtime="00:03:04.18" resultid="4159" heatid="6280" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:29.26" />
                    <SPLIT distance="150" swimtime="00:02:17.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="698" reactiontime="+82" swimtime="00:00:33.98" resultid="4160" heatid="6345" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1610" points="842" reactiontime="+96" swimtime="00:01:32.68" resultid="4161" heatid="6400" lane="2" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="STANISŁAW" gender="M" lastname="KISZCZAK" nation="POL" athleteid="4162">
              <RESULTS>
                <RESULT eventid="1528" points="566" reactiontime="+105" swimtime="00:00:32.99" resultid="4163" heatid="6346" lane="1" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="GRAŻYNA" gender="F" lastname="KISZCZAK" nation="POL" athleteid="4164">
              <RESULTS>
                <RESULT eventid="1153" points="848" reactiontime="+82" swimtime="00:01:26.64" resultid="4165" heatid="6078" lane="3" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. H" eventid="1213" points="1007" reactiontime="+75" swimtime="00:00:38.33" resultid="4166" heatid="6123" lane="4" entrytime="00:00:40.00" />
                <RESULT comment="Rekord Polski kat. H" eventid="1348" points="805" reactiontime="+82" swimtime="00:00:39.32" resultid="4167" heatid="6220" lane="1" entrytime="00:00:40.00" />
                <RESULT comment="Rekord Polski kat. H" eventid="1452" points="739" reactiontime="+84" swimtime="00:03:19.37" resultid="4168" heatid="6295" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.56" />
                    <SPLIT distance="100" swimtime="00:01:36.52" />
                    <SPLIT distance="150" swimtime="00:02:32.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="776" reactiontime="+81" swimtime="00:00:34.98" resultid="4169" heatid="6335" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1543" points="906" reactiontime="+81" swimtime="00:03:15.46" resultid="4170" heatid="6370" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                    <SPLIT distance="100" swimtime="00:01:36.58" />
                    <SPLIT distance="150" swimtime="00:02:27.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-01" firstname="RENATA" gender="F" lastname="BASTEK" nation="POL" athleteid="4171">
              <RESULTS>
                <RESULT eventid="1213" points="851" reactiontime="+67" swimtime="00:00:43.41" resultid="4172" heatid="6122" lane="5" entrytime="00:00:44.00" />
                <RESULT eventid="1348" points="642" reactiontime="+76" swimtime="00:00:45.49" resultid="4173" heatid="6219" lane="4" entrytime="00:00:46.00" />
                <RESULT eventid="1513" points="963" reactiontime="+78" swimtime="00:00:35.22" resultid="4174" heatid="6334" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-01" firstname="KRYSTYNA" gender="F" lastname="FECICA" nation="POL" athleteid="4175">
              <RESULTS>
                <RESULT eventid="1183" points="741" reactiontime="+105" swimtime="00:03:59.06" resultid="4176" heatid="6104" lane="2" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.69" />
                    <SPLIT distance="100" swimtime="00:01:55.80" />
                    <SPLIT distance="150" swimtime="00:02:58.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="630" reactiontime="+104" swimtime="00:00:51.13" resultid="4177" heatid="6196" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1483" points="479" swimtime="00:01:50.46" resultid="4178" heatid="6313" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="640" reactiontime="+100" swimtime="00:01:52.77" resultid="4179" heatid="6505" lane="3" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-01-01" firstname="DANIEL" gender="M" lastname="FECICA" nation="POL" athleteid="4180">
              <RESULTS>
                <RESULT eventid="1198" points="808" reactiontime="+99" swimtime="00:03:29.28" resultid="4181" heatid="6111" lane="5" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                    <SPLIT distance="100" swimtime="00:01:42.14" />
                    <SPLIT distance="150" swimtime="00:02:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="642" reactiontime="+92" swimtime="00:00:44.30" resultid="4182" heatid="6208" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="1610" points="741" reactiontime="+97" swimtime="00:01:36.72" resultid="4183" heatid="6399" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="BERNARD" gender="M" lastname="POLOCZEK" nation="POL" athleteid="4184">
              <RESULTS>
                <RESULT eventid="1228" points="609" reactiontime="+62" swimtime="00:00:41.62" resultid="4185" heatid="6130" lane="2" entrytime="00:00:42.01" />
                <RESULT eventid="1393" points="615" reactiontime="+58" swimtime="00:01:34.01" resultid="4186" heatid="6253" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="539" reactiontime="+65" swimtime="00:03:34.47" resultid="4187" heatid="6374" lane="5" entrytime="00:03:42.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.15" />
                    <SPLIT distance="100" swimtime="00:01:41.32" />
                    <SPLIT distance="150" swimtime="00:02:38.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="BARBARA" gender="F" lastname="BRENDLER" nation="POL" athleteid="4188">
              <RESULTS>
                <RESULT eventid="1153" points="307" reactiontime="+103" swimtime="00:02:01.50" resultid="4189" heatid="6075" lane="4" entrytime="00:01:56.00" />
                <RESULT eventid="1257" points="482" reactiontime="+98" swimtime="00:01:31.05" resultid="4190" heatid="6150" lane="3" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="445" reactiontime="+78" swimtime="00:03:32.12" resultid="4191" heatid="6272" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                    <SPLIT distance="100" swimtime="00:01:39.07" />
                    <SPLIT distance="150" swimtime="00:02:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="516" reactiontime="+92" swimtime="00:00:40.06" resultid="4192" heatid="6332" lane="5" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="BEATA" gender="F" lastname="SULEWSKA" nation="POL" athleteid="4193">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. D" eventid="1058" points="776" reactiontime="+96" swimtime="00:05:46.25" resultid="4194" heatid="6431" lane="2" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                    <SPLIT distance="100" swimtime="00:01:18.76" />
                    <SPLIT distance="150" swimtime="00:02:06.34" />
                    <SPLIT distance="200" swimtime="00:02:52.79" />
                    <SPLIT distance="250" swimtime="00:03:39.89" />
                    <SPLIT distance="300" swimtime="00:04:28.99" />
                    <SPLIT distance="350" swimtime="00:05:07.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="727" reactiontime="+99" swimtime="00:03:01.56" resultid="4195" heatid="6107" lane="5" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.20" />
                    <SPLIT distance="100" swimtime="00:01:28.35" />
                    <SPLIT distance="150" swimtime="00:02:14.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="613" reactiontime="+92" swimtime="00:01:09.41" resultid="4196" heatid="6157" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="4197" heatid="6200" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1452" points="707" reactiontime="+96" swimtime="00:02:45.84" resultid="4198" heatid="6298" lane="1" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:01:21.17" />
                    <SPLIT distance="150" swimtime="00:02:07.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="634" reactiontime="+93" swimtime="00:01:27.46" resultid="4199" heatid="6510" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="700" reactiontime="+88" swimtime="00:05:06.33" resultid="4200" heatid="6558" lane="4" entrytime="00:05:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:01:13.05" />
                    <SPLIT distance="150" swimtime="00:01:51.98" />
                    <SPLIT distance="200" swimtime="00:02:31.40" />
                    <SPLIT distance="250" swimtime="00:03:10.67" />
                    <SPLIT distance="300" swimtime="00:03:50.16" />
                    <SPLIT distance="350" swimtime="00:04:29.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="MAREK" gender="M" lastname="ROTHER" nation="POL" athleteid="4201">
              <RESULTS>
                <RESULT eventid="1228" points="783" reactiontime="+64" swimtime="00:00:30.40" resultid="4202" heatid="6137" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="1272" points="635" reactiontime="+86" swimtime="00:01:02.12" resultid="4203" heatid="6172" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="793" reactiontime="+63" swimtime="00:01:05.59" resultid="4204" heatid="6261" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="641" reactiontime="+86" swimtime="00:02:17.26" resultid="4205" heatid="6289" lane="5" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:06.67" />
                    <SPLIT distance="150" swimtime="00:01:41.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="797" reactiontime="+60" swimtime="00:02:26.14" resultid="4206" heatid="6382" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:49.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="MARTA" gender="F" lastname="FRANK" nation="POL" athleteid="4207">
              <RESULTS>
                <RESULT eventid="1153" points="598" reactiontime="+79" swimtime="00:01:21.12" resultid="4208" heatid="6081" lane="5" entrytime="00:01:19.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="646" reactiontime="+63" swimtime="00:00:36.35" resultid="4209" heatid="6124" lane="4" entrytime="00:00:36.29" />
                <RESULT eventid="1378" points="552" reactiontime="+68" swimtime="00:01:21.25" resultid="4210" heatid="6247" lane="4" entrytime="00:01:20.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="501" reactiontime="+82" swimtime="00:03:06.07" resultid="4211" heatid="6297" lane="5" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:26.74" />
                    <SPLIT distance="150" swimtime="00:02:21.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="558" reactiontime="+76" swimtime="00:00:33.02" resultid="4212" heatid="6338" lane="5" entrytime="00:00:31.01" />
                <RESULT eventid="1543" points="512" reactiontime="+73" swimtime="00:03:01.78" resultid="4213" heatid="6370" lane="4" entrytime="00:03:04.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:01:28.23" />
                    <SPLIT distance="150" swimtime="00:02:15.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="WŁODZIMIERZ" gender="M" lastname="BOSOWSKI" nation="POL" athleteid="4214">
              <RESULTS>
                <RESULT eventid="1168" points="310" reactiontime="+98" swimtime="00:01:46.16" resultid="4215" heatid="6085" lane="1" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="244" reactiontime="+94" swimtime="00:00:53.50" resultid="4216" heatid="6128" lane="3" entrytime="00:00:48.50" />
                <RESULT eventid="1363" points="410" reactiontime="+106" swimtime="00:00:40.85" resultid="4217" heatid="6226" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1528" points="396" reactiontime="+91" swimtime="00:00:37.16" resultid="4218" heatid="6344" lane="5" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="JANINA" gender="F" lastname="BOSOWSKA" nation="POL" athleteid="4219">
              <RESULTS>
                <RESULT eventid="1153" points="522" reactiontime="+86" swimtime="00:01:52.88" resultid="4220" heatid="6075" lane="5" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="513" reactiontime="+62" swimtime="00:00:51.36" resultid="4221" heatid="6120" lane="6" entrytime="00:00:58.00" />
                <RESULT eventid="1318" points="630" reactiontime="+83" swimtime="00:00:51.14" resultid="4222" heatid="6195" lane="3" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="WIESŁAW" gender="M" lastname="KORNICKI" nation="POL" athleteid="4223">
              <RESULTS>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="4224" heatid="6347" lane="4" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="MARTA" gender="F" lastname="ORACZ" nation="POL" athleteid="4225">
              <RESULTS>
                <RESULT eventid="1122" points="315" swimtime="00:13:51.34" resultid="4226" heatid="6442" lane="3" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                    <SPLIT distance="100" swimtime="00:01:31.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="DOROTA" gender="F" lastname="KRAUZE" nation="POL" athleteid="4227">
              <RESULTS>
                <RESULT eventid="1183" status="DNS" swimtime="00:00:00.00" resultid="4228" heatid="6103" lane="1" entrytime="00:04:35.00" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="4229" heatid="6195" lane="5" entrytime="00:00:53.00" />
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="4230" heatid="6505" lane="2" entrytime="00:01:59.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="MACIEJ" gender="M" lastname="KUNICKI" nation="POL" athleteid="4231">
              <RESULTS>
                <RESULT eventid="1302" points="451" reactiontime="+88" swimtime="00:02:50.04" resultid="4232" heatid="6189" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:20.18" />
                    <SPLIT distance="150" swimtime="00:02:06.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="615" reactiontime="+89" swimtime="00:00:31.35" resultid="4233" heatid="6235" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1498" points="570" reactiontime="+93" swimtime="00:01:10.72" resultid="4234" heatid="6322" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="ALEKSANDRA" gender="F" lastname="TUSZYŃSKA" nation="POL" athleteid="4235">
              <RESULTS>
                <RESULT eventid="1213" points="581" reactiontime="+71" swimtime="00:00:37.51" resultid="4236" heatid="6124" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1257" points="511" reactiontime="+100" swimtime="00:01:12.17" resultid="4237" heatid="6157" lane="6" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="618" reactiontime="+91" swimtime="00:00:34.32" resultid="4238" heatid="6222" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1513" points="658" reactiontime="+92" swimtime="00:00:30.81" resultid="4239" heatid="6339" lane="2" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="RYSZARD" gender="M" lastname="TYLEK" nation="POL" athleteid="4240">
              <RESULTS>
                <RESULT eventid="1333" points="362" reactiontime="+101" swimtime="00:00:48.04" resultid="4241" heatid="6209" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1610" status="DNS" swimtime="00:00:00.00" resultid="4242" heatid="6397" lane="4" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="DANIEL" gender="M" lastname="WESELAK" nation="POL" athleteid="4243">
              <RESULTS>
                <RESULT eventid="1168" points="489" reactiontime="+86" swimtime="00:01:13.95" resultid="4244" heatid="6094" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" status="DNS" swimtime="00:00:00.00" resultid="4245" heatid="6235" lane="3" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="DANIEL" gender="M" lastname="HOSZCZEWSKI" nation="POL" athleteid="4246">
              <RESULTS>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="4247" heatid="6175" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="1363" status="DNS" swimtime="00:00:00.00" resultid="4248" heatid="6235" lane="2" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+60" swimtime="00:02:47.09" resultid="4253" heatid="6522" lane="3" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                    <SPLIT distance="100" swimtime="00:01:30.28" />
                    <SPLIT distance="150" swimtime="00:02:13.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4184" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="4240" number="2" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4214" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4162" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+81" swimtime="00:02:32.13" resultid="4254" heatid="6523" lane="5" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                    <SPLIT distance="100" swimtime="00:01:28.86" />
                    <SPLIT distance="150" swimtime="00:01:59.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4155" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4180" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4231" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4139" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+87" swimtime="00:02:14.11" resultid="4257" heatid="6532" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:45.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4223" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="4155" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4162" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="4201" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="10">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+100" swimtime="00:02:16.31" resultid="4258" heatid="6531" lane="5" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:01:42.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4214" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="4184" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="4231" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4139" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1243" reactiontime="+63" swimtime="00:02:49.91" resultid="4251" heatid="6519" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.04" />
                    <SPLIT distance="150" swimtime="00:02:11.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4171" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4151" number="2" />
                    <RELAYPOSITION athleteid="4164" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="4188" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="1243" reactiontime="+81" swimtime="00:02:30.09" resultid="4252" heatid="6520" lane="2" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                    <SPLIT distance="100" swimtime="00:01:23.84" />
                    <SPLIT distance="150" swimtime="00:01:58.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4146" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4193" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="4235" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4207" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="7">
              <RESULTS>
                <RESULT eventid="1408" swimtime="00:02:39.02" resultid="4255" heatid="6527" lane="2" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                    <SPLIT distance="100" swimtime="00:01:27.01" />
                    <SPLIT distance="150" swimtime="00:02:02.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4188" number="1" />
                    <RELAYPOSITION athleteid="4175" number="2" />
                    <RELAYPOSITION athleteid="4171" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="4164" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="8">
              <RESULTS>
                <RESULT eventid="1408" reactiontime="+89" swimtime="00:02:14.80" resultid="4256" heatid="6528" lane="4" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:11.13" />
                    <SPLIT distance="150" swimtime="00:01:44.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4146" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="4193" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="4207" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="4235" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+93" swimtime="00:02:33.30" resultid="4249" heatid="6495" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.18" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                    <SPLIT distance="150" swimtime="00:01:57.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4219" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="4146" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="4214" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="4223" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+92" swimtime="00:02:19.38" resultid="4250" heatid="6496" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:16.30" />
                    <SPLIT distance="150" swimtime="00:01:47.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4188" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="4184" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4235" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="4139" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="11">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+70" swimtime="00:02:50.27" resultid="4259" heatid="6535" lane="3" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:01:27.12" />
                    <SPLIT distance="150" swimtime="00:02:16.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4171" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4180" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="4175" number="3" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4155" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="12">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+76" swimtime="00:02:40.12" resultid="4260" heatid="6536" lane="3" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:26.75" />
                    <SPLIT distance="150" swimtime="00:02:07.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4164" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4151" number="2" reactiontime="+85" />
                    <RELAYPOSITION athleteid="4214" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="4139" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="13">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+74" swimtime="00:02:13.62" resultid="4261" heatid="6538" lane="3" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:12.34" />
                    <SPLIT distance="150" swimtime="00:01:43.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4201" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4207" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4231" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="4235" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WMT" name="Warsaw Masters Team" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" email="jstobnic@gmail.com" name="Justyna Marta Stobnicka" state="MAZ" />
          <ATHLETES>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="4289">
              <RESULTS>
                <RESULT eventid="1092" points="400" reactiontime="+112" swimtime="00:09:19.76" resultid="4290" heatid="6486" lane="1" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.21" />
                    <SPLIT distance="100" swimtime="00:02:21.06" />
                    <SPLIT distance="150" swimtime="00:03:35.27" />
                    <SPLIT distance="200" swimtime="00:04:48.39" />
                    <SPLIT distance="250" swimtime="00:05:57.89" />
                    <SPLIT distance="300" swimtime="00:07:11.28" />
                    <SPLIT distance="350" swimtime="00:08:14.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="384" reactiontime="+116" swimtime="00:04:37.05" resultid="4291" heatid="6109" lane="1" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.33" />
                    <SPLIT distance="100" swimtime="00:02:14.88" />
                    <SPLIT distance="150" swimtime="00:03:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="281" reactiontime="+123" swimtime="00:05:15.59" resultid="4292" heatid="6183" lane="4" entrytime="00:05:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.51" />
                    <SPLIT distance="100" swimtime="00:02:33.19" />
                    <SPLIT distance="150" swimtime="00:03:56.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="430" reactiontime="+117" swimtime="00:00:53.11" resultid="4293" heatid="6203" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="1467" points="357" reactiontime="+117" swimtime="00:04:27.73" resultid="4294" heatid="6299" lane="4" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.76" />
                    <SPLIT distance="100" swimtime="00:02:10.57" />
                    <SPLIT distance="150" swimtime="00:03:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="240" reactiontime="+119" swimtime="00:02:27.97" resultid="4295" heatid="6316" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="389" reactiontime="+119" swimtime="00:02:01.35" resultid="4296" heatid="6395" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-28" firstname="Monika" gender="F" lastname="Figura" nation="POL" athleteid="4297">
              <RESULTS>
                <RESULT eventid="1122" status="DNS" swimtime="00:00:00.00" resultid="4298" heatid="6444" lane="3" entrytime="00:11:58.00" />
                <RESULT eventid="1213" points="598" reactiontime="+78" swimtime="00:00:37.15" resultid="4299" heatid="6124" lane="5" entrytime="00:00:37.12" />
                <RESULT eventid="1257" points="509" reactiontime="+75" swimtime="00:01:12.29" resultid="4300" heatid="6155" lane="3" entrytime="00:01:13.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="463" reactiontime="+80" swimtime="00:01:23.67" resultid="4301" heatid="6247" lane="5" entrytime="00:01:22.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="4302" heatid="6276" lane="6" entrytime="00:02:49.76" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="4303" heatid="6369" lane="2" entrytime="00:03:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="4304">
              <RESULTS>
                <RESULT eventid="1168" points="933" reactiontime="+77" swimtime="00:01:07.05" resultid="4305" heatid="6097" lane="5" entrytime="00:01:07.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="967" reactiontime="+77" swimtime="00:00:57.53" resultid="4306" heatid="6178" lane="1" entrytime="00:00:57.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="792" reactiontime="+77" swimtime="00:00:29.97" resultid="4307" heatid="6237" lane="5" entrytime="00:00:29.83" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="4308" heatid="6290" lane="6" entrytime="00:02:12.11" />
                <RESULT eventid="1528" points="842" reactiontime="+78" swimtime="00:00:26.86" resultid="4309" heatid="6360" lane="4" entrytime="00:00:26.85" />
                <RESULT eventid="1610" status="DNS" swimtime="00:00:00.00" resultid="4310" heatid="6406" lane="1" entrytime="00:01:17.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-02" firstname="Maciej" gender="M" lastname="Falkowski" nation="POL" athleteid="4311">
              <RESULTS>
                <RESULT eventid="1168" points="657" reactiontime="+86" swimtime="00:01:06.59" resultid="4312" heatid="6097" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="701" reactiontime="+83" swimtime="00:00:56.93" resultid="4313" heatid="6178" lane="2" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="742" reactiontime="+83" swimtime="00:00:28.01" resultid="4314" heatid="6233" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1528" points="696" reactiontime="+83" swimtime="00:00:25.65" resultid="4315" heatid="6361" lane="4" entrytime="00:00:26.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="4316">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. C" eventid="1228" points="1078" reactiontime="+66" swimtime="00:00:26.80" resultid="4317" heatid="6139" lane="5" entrytime="00:00:27.99" />
                <RESULT eventid="1363" points="873" reactiontime="+80" swimtime="00:00:26.30" resultid="4318" heatid="6241" lane="4" entrytime="00:00:26.49" />
                <RESULT comment="Rekord Polski kat. C" eventid="1393" points="916" reactiontime="+65" swimtime="00:01:00.54" resultid="4319" heatid="6262" lane="5" entrytime="00:01:01.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="4320" heatid="6327" lane="6" entrytime="00:00:59.59" />
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="4321" heatid="6382" lane="1" entrytime="00:02:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-07-15" firstname="Piotr" gender="M" lastname="Kober" nation="POL" athleteid="4322">
              <RESULTS>
                <RESULT eventid="1137" points="215" swimtime="00:14:23.44" resultid="4323" heatid="6448" lane="1" entrytime="00:14:47.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.50" />
                    <SPLIT distance="100" swimtime="00:01:42.37" />
                    <SPLIT distance="200" swimtime="00:03:33.82" />
                    <SPLIT distance="300" swimtime="00:05:24.56" />
                    <SPLIT distance="400" swimtime="00:07:15.35" />
                    <SPLIT distance="500" swimtime="00:09:02.65" />
                    <SPLIT distance="600" swimtime="00:10:48.56" />
                    <SPLIT distance="700" swimtime="00:12:38.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="214" reactiontime="+130" swimtime="00:01:43.12" resultid="4324" heatid="6085" lane="6" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="183" reactiontime="+116" swimtime="00:00:49.28" resultid="4325" heatid="6129" lane="1" entrytime="00:00:46.41" />
                <RESULT eventid="1333" points="176" reactiontime="+86" swimtime="00:00:52.60" resultid="4326" heatid="6203" lane="1" entrytime="00:00:56.78" />
                <RESULT eventid="1437" points="211" reactiontime="+107" swimtime="00:03:18.81" resultid="4327" heatid="6279" lane="5" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                    <SPLIT distance="100" swimtime="00:01:35.16" />
                    <SPLIT distance="150" swimtime="00:02:28.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="4328" heatid="6343" lane="5" entrytime="00:00:41.12" />
                <RESULT eventid="1640" status="DNS" swimtime="00:00:00.00" resultid="4329" heatid="6561" lane="5" entrytime="00:07:00.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="4330">
              <RESULTS>
                <RESULT eventid="1168" points="809" reactiontime="+85" swimtime="00:01:08.25" resultid="4331" heatid="6098" lane="6" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="814" reactiontime="+76" swimtime="00:00:30.90" resultid="4332" heatid="6136" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1393" points="865" reactiontime="+74" swimtime="00:01:08.28" resultid="4333" heatid="6261" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="777" reactiontime="+90" swimtime="00:02:32.06" resultid="4334" heatid="6309" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:10.12" />
                    <SPLIT distance="150" swimtime="00:01:56.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="696" reactiontime="+84" swimtime="00:00:27.67" resultid="4335" heatid="6348" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1558" points="806" reactiontime="+80" swimtime="00:02:31.42" resultid="4336" heatid="6380" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:14.47" />
                    <SPLIT distance="150" swimtime="00:01:53.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="4337">
              <RESULTS>
                <RESULT eventid="1198" points="399" reactiontime="+102" swimtime="00:03:29.02" resultid="4338" heatid="6112" lane="6" entrytime="00:03:24.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.72" />
                    <SPLIT distance="100" swimtime="00:01:38.12" />
                    <SPLIT distance="150" swimtime="00:02:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="149" reactiontime="+104" swimtime="00:00:54.36" resultid="4339" heatid="6127" lane="3" entrytime="00:00:53.74" />
                <RESULT eventid="1333" points="375" swimtime="00:00:42.57" resultid="4340" heatid="6206" lane="2" entrytime="00:00:44.26" />
                <RESULT eventid="1393" points="143" reactiontime="+118" swimtime="00:02:04.36" resultid="4341" heatid="6251" lane="5" entrytime="00:01:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="258" reactiontime="+101" swimtime="00:00:38.50" resultid="4342" heatid="6344" lane="1" entrytime="00:00:37.26" />
                <RESULT eventid="1610" points="388" reactiontime="+96" swimtime="00:01:34.22" resultid="4343" heatid="6398" lane="2" entrytime="00:01:37.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-05-05" firstname="Dominik" gender="M" lastname="Matuzewicz" nation="POL" athleteid="4344">
              <RESULTS>
                <RESULT eventid="1528" points="723" reactiontime="+79" swimtime="00:00:25.70" resultid="4345" heatid="6364" lane="6" entrytime="00:00:25.86" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-29" firstname="Jan Maciej" gender="M" lastname="Boboli" nation="POL" athleteid="4346">
              <RESULTS>
                <RESULT eventid="1228" points="173" reactiontime="+82" swimtime="00:00:59.97" resultid="4347" heatid="6127" lane="2" entrytime="00:00:56.00" />
                <RESULT eventid="1272" points="285" reactiontime="+103" swimtime="00:01:34.75" resultid="4348" heatid="6161" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="430" reactiontime="+115" swimtime="00:00:40.21" resultid="4349" heatid="6226" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1437" points="203" reactiontime="+106" swimtime="00:03:59.93" resultid="4350" heatid="6280" lane="4" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                    <SPLIT distance="100" swimtime="00:01:45.41" />
                    <SPLIT distance="150" swimtime="00:02:52.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="419" reactiontime="+99" swimtime="00:00:36.46" resultid="4351" heatid="6346" lane="5" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-14" firstname="Wojciech" gender="M" lastname="Kałużyński" nation="POL" athleteid="4352">
              <RESULTS>
                <RESULT eventid="1137" points="372" swimtime="00:11:33.02" resultid="4353" heatid="6453" lane="4" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.20" />
                    <SPLIT distance="200" swimtime="00:02:43.90" />
                    <SPLIT distance="300" swimtime="00:04:13.61" />
                    <SPLIT distance="400" swimtime="00:05:45.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="381" reactiontime="+87" swimtime="00:01:20.32" resultid="4354" heatid="6089" lane="4" entrytime="00:01:21.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="420" reactiontime="+83" swimtime="00:01:07.61" resultid="4355" heatid="6168" lane="3" entrytime="00:01:07.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="364" reactiontime="+84" swimtime="00:02:36.25" resultid="4356" heatid="6284" lane="3" entrytime="00:02:34.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                    <SPLIT distance="150" swimtime="00:01:54.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="462" reactiontime="+83" swimtime="00:00:29.83" resultid="4357" heatid="6352" lane="6" entrytime="00:00:30.10" />
                <RESULT eventid="1640" points="374" reactiontime="+86" swimtime="00:05:33.93" resultid="4358" heatid="6565" lane="1" entrytime="00:05:36.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                    <SPLIT distance="150" swimtime="00:02:02.16" />
                    <SPLIT distance="200" swimtime="00:02:44.60" />
                    <SPLIT distance="250" swimtime="00:04:10.51" />
                    <SPLIT distance="300" swimtime="00:04:53.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-12-31" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="4359">
              <RESULTS>
                <RESULT eventid="1168" points="818" reactiontime="+88" swimtime="00:01:12.73" resultid="4360" heatid="6092" lane="3" entrytime="00:01:14.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="832" reactiontime="+89" swimtime="00:01:02.39" resultid="4361" heatid="6171" lane="6" entrytime="00:01:04.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="743" reactiontime="+81" swimtime="00:01:14.59" resultid="4362" heatid="6256" lane="3" entrytime="00:01:17.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="883" reactiontime="+85" swimtime="00:02:41.31" resultid="4363" heatid="6307" lane="4" entrytime="00:02:41.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:02:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="806" reactiontime="+75" swimtime="00:02:41.79" resultid="4364" heatid="6380" lane="1" entrytime="00:02:39.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                    <SPLIT distance="100" swimtime="00:01:18.59" />
                    <SPLIT distance="150" swimtime="00:02:00.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="Borodziuk" nation="POL" athleteid="4365">
              <RESULTS>
                <RESULT eventid="1137" points="369" swimtime="00:15:46.72" resultid="4366" heatid="6448" lane="6" entrytime="00:15:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                    <SPLIT distance="100" swimtime="00:01:42.68" />
                    <SPLIT distance="200" swimtime="00:03:37.74" />
                    <SPLIT distance="300" swimtime="00:05:37.57" />
                    <SPLIT distance="400" swimtime="00:07:40.84" />
                    <SPLIT distance="500" swimtime="00:09:45.01" />
                    <SPLIT distance="600" swimtime="00:11:49.83" />
                    <SPLIT distance="700" swimtime="00:13:52.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="432" reactiontime="+84" swimtime="00:00:46.67" resultid="4367" heatid="6129" lane="6" entrytime="00:00:47.00" />
                <RESULT eventid="1272" points="508" reactiontime="+93" swimtime="00:01:22.74" resultid="4368" heatid="6161" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="322" reactiontime="+84" swimtime="00:00:52.79" resultid="4369" heatid="6203" lane="3" entrytime="00:00:54.00" />
                <RESULT eventid="1437" points="468" reactiontime="+100" swimtime="00:03:11.42" resultid="4370" heatid="6280" lane="1" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:32.02" />
                    <SPLIT distance="150" swimtime="00:02:22.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="4371" heatid="6344" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1640" points="417" reactiontime="+94" swimtime="00:07:17.76" resultid="4372" heatid="6561" lane="1" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.82" />
                    <SPLIT distance="100" swimtime="00:01:38.03" />
                    <SPLIT distance="150" swimtime="00:02:34.70" />
                    <SPLIT distance="200" swimtime="00:03:31.95" />
                    <SPLIT distance="250" swimtime="00:04:29.98" />
                    <SPLIT distance="300" swimtime="00:05:28.26" />
                    <SPLIT distance="350" swimtime="00:06:25.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-12-31" firstname="Paweł" gender="M" lastname="Kowalewski" nation="POL" athleteid="4373">
              <RESULTS>
                <RESULT eventid="1467" points="830" reactiontime="+79" swimtime="00:02:28.76" resultid="6551" heatid="6311" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="150" swimtime="00:01:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat.E" eventid="1137" points="824" swimtime="00:09:46.80" resultid="4374" heatid="6454" lane="3" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="200" swimtime="00:02:19.46" />
                    <SPLIT distance="300" swimtime="00:03:31.80" />
                    <SPLIT distance="400" swimtime="00:05:59.97" />
                    <SPLIT distance="500" swimtime="00:05:59.97" />
                    <SPLIT distance="600" swimtime="00:07:14.62" />
                    <SPLIT distance="700" swimtime="00:08:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. E" eventid="1437" points="845" reactiontime="+77" swimtime="00:02:09.61" resultid="4375" heatid="6281" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                    <SPLIT distance="100" swimtime="00:01:03.21" />
                    <SPLIT distance="150" swimtime="00:01:36.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="703" reactiontime="+77" swimtime="00:01:08.96" resultid="4377" heatid="6323" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="838" reactiontime="+74" swimtime="00:04:38.70" resultid="4378" heatid="6568" lane="5" entrytime="00:04:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:05.93" />
                    <SPLIT distance="150" swimtime="00:01:41.43" />
                    <SPLIT distance="200" swimtime="00:02:16.90" />
                    <SPLIT distance="250" swimtime="00:02:52.14" />
                    <SPLIT distance="300" swimtime="00:03:27.19" />
                    <SPLIT distance="350" swimtime="00:04:02.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="4379">
              <RESULTS>
                <RESULT eventid="1183" points="717" reactiontime="+96" swimtime="00:03:11.26" resultid="4380" heatid="6107" lane="1" entrytime="00:03:06.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="100" swimtime="00:01:31.26" />
                    <SPLIT distance="150" swimtime="00:02:21.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="591" reactiontime="+89" swimtime="00:01:15.69" resultid="4381" heatid="6155" lane="2" entrytime="00:01:13.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="700" reactiontime="+85" swimtime="00:00:40.62" resultid="4382" heatid="6200" lane="4" entrytime="00:00:39.43" />
                <RESULT eventid="1422" points="561" reactiontime="+87" swimtime="00:02:47.26" resultid="4383" heatid="6276" lane="5" entrytime="00:02:41.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                    <SPLIT distance="100" swimtime="00:01:21.87" />
                    <SPLIT distance="150" swimtime="00:02:06.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="552" reactiontime="+83" swimtime="00:00:34.32" resultid="4384" heatid="6336" lane="5" entrytime="00:00:34.08" />
                <RESULT eventid="1595" points="744" reactiontime="+82" swimtime="00:01:27.47" resultid="4385" heatid="6509" lane="3" entrytime="00:01:26.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-12-31" firstname="Robert" gender="M" lastname="Nowicki" nation="POL" athleteid="4386">
              <RESULTS>
                <RESULT eventid="1272" points="222" reactiontime="+100" swimtime="00:01:30.45" resultid="4387" heatid="6160" lane="4" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-12-31" firstname="Katarzyna" gender="F" lastname="Dobczyńska" nation="POL" athleteid="4388">
              <RESULTS>
                <RESULT eventid="1213" points="363" reactiontime="+81" swimtime="00:00:43.88" resultid="4389" heatid="6121" lane="2" entrytime="00:00:46.00" />
                <RESULT eventid="1257" points="327" reactiontime="+100" swimtime="00:01:23.73" resultid="4390" heatid="6152" lane="6" entrytime="00:01:26.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" status="DNS" swimtime="00:00:00.00" resultid="4391" heatid="6246" lane="2" entrytime="00:01:33.08" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-12-31" firstname="Arkadiusz" gender="M" lastname="Dobrzyński" nation="POL" athleteid="4392">
              <RESULTS>
                <RESULT eventid="1228" points="621" reactiontime="+72" swimtime="00:00:32.21" resultid="4393" heatid="6136" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="4394" heatid="6173" lane="4" entrytime="00:01:01.00" />
                <RESULT eventid="1363" points="541" reactiontime="+82" swimtime="00:00:30.84" resultid="4395" heatid="6234" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1393" points="603" reactiontime="+74" swimtime="00:01:09.59" resultid="4396" heatid="6260" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="590" reactiontime="+73" swimtime="00:00:27.59" resultid="4397" heatid="6361" lane="5" entrytime="00:00:26.70" />
                <RESULT eventid="1558" points="517" reactiontime="+75" swimtime="00:02:38.39" resultid="4398" heatid="6379" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:17.91" />
                    <SPLIT distance="150" swimtime="00:01:58.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-06-16" firstname="Elżbieta" gender="F" lastname="Janik" nation="POL" athleteid="4399">
              <RESULTS>
                <RESULT eventid="1378" points="416" reactiontime="+77" swimtime="00:02:23.61" resultid="4400" heatid="6243" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="149" reactiontime="+112" swimtime="00:01:15.92" resultid="4401" heatid="6328" lane="3" entrytime="00:01:18.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-06-02" firstname="Wojciech" gender="M" lastname="Czupryn" nation="POL" athleteid="4402">
              <RESULTS>
                <RESULT eventid="1137" points="323" swimtime="00:13:45.97" resultid="4403" heatid="6449" lane="1" entrytime="00:13:52.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                    <SPLIT distance="100" swimtime="00:01:39.10" />
                    <SPLIT distance="200" swimtime="00:03:23.16" />
                    <SPLIT distance="300" swimtime="00:05:07.00" />
                    <SPLIT distance="400" swimtime="00:06:51.58" />
                    <SPLIT distance="500" swimtime="00:10:20.86" />
                    <SPLIT distance="600" swimtime="00:10:20.86" />
                    <SPLIT distance="700" swimtime="00:12:04.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="319" reactiontime="+92" swimtime="00:01:35.83" resultid="4404" heatid="6085" lane="3" entrytime="00:01:37.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="358" reactiontime="+90" swimtime="00:01:20.08" resultid="4405" heatid="6162" lane="2" entrytime="00:01:17.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="327" reactiontime="+97" swimtime="00:00:46.70" resultid="4406" heatid="6205" lane="6" entrytime="00:00:47.63" />
                <RESULT eventid="1393" points="258" reactiontime="+89" swimtime="00:01:45.44" resultid="4407" heatid="6251" lane="1" entrytime="00:01:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="284" reactiontime="+86" swimtime="00:03:46.52" resultid="4408" heatid="6373" lane="2" entrytime="00:04:05.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.82" />
                    <SPLIT distance="100" swimtime="00:01:51.91" />
                    <SPLIT distance="150" swimtime="00:02:50.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="342" reactiontime="+104" swimtime="00:06:23.68" resultid="4409" heatid="6562" lane="2" entrytime="00:06:21.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="150" swimtime="00:02:20.78" />
                    <SPLIT distance="200" swimtime="00:03:10.54" />
                    <SPLIT distance="250" swimtime="00:04:00.01" />
                    <SPLIT distance="300" swimtime="00:04:49.29" />
                    <SPLIT distance="350" swimtime="00:05:38.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-13" firstname="Ewa" gender="F" lastname="Krzyżanowska" nation="POL" athleteid="4410">
              <RESULTS>
                <RESULT eventid="1122" points="360" swimtime="00:13:15.14" resultid="4411" heatid="6443" lane="3" entrytime="00:13:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:30.24" />
                    <SPLIT distance="200" swimtime="00:03:09.50" />
                    <SPLIT distance="300" swimtime="00:04:49.99" />
                    <SPLIT distance="400" swimtime="00:06:32.61" />
                    <SPLIT distance="500" swimtime="00:08:15.99" />
                    <SPLIT distance="600" swimtime="00:09:56.98" />
                    <SPLIT distance="700" swimtime="00:11:38.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="516" reactiontime="+80" swimtime="00:00:39.18" resultid="4412" heatid="6123" lane="5" entrytime="00:00:40.55" />
                <RESULT eventid="1257" points="512" reactiontime="+97" swimtime="00:01:13.68" resultid="4413" heatid="6154" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="442" reactiontime="+93" swimtime="00:02:50.52" resultid="4414" heatid="6275" lane="6" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:21.61" />
                    <SPLIT distance="150" swimtime="00:02:06.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="579" reactiontime="+91" swimtime="00:00:32.62" resultid="4415" heatid="6337" lane="1" entrytime="00:00:33.08" />
                <RESULT eventid="1625" points="371" reactiontime="+97" swimtime="00:06:18.39" resultid="4416" heatid="6556" lane="1" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                    <SPLIT distance="100" swimtime="00:01:26.08" />
                    <SPLIT distance="150" swimtime="00:02:14.60" />
                    <SPLIT distance="200" swimtime="00:03:03.82" />
                    <SPLIT distance="250" swimtime="00:03:53.58" />
                    <SPLIT distance="300" swimtime="00:04:42.86" />
                    <SPLIT distance="350" swimtime="00:05:31.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-12-31" firstname="Anna" gender="F" lastname="Stanisławska" nation="POL" athleteid="4417">
              <RESULTS>
                <RESULT eventid="1058" points="253" reactiontime="+112" swimtime="00:07:58.66" resultid="4418" heatid="6428" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="100" swimtime="00:01:46.32" />
                    <SPLIT distance="150" swimtime="00:02:51.30" />
                    <SPLIT distance="200" swimtime="00:03:56.82" />
                    <SPLIT distance="250" swimtime="00:05:03.54" />
                    <SPLIT distance="300" swimtime="00:06:08.41" />
                    <SPLIT distance="350" swimtime="00:07:04.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="258" reactiontime="+90" swimtime="00:01:42.95" resultid="4419" heatid="6077" lane="1" entrytime="00:01:41.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="288" reactiontime="+93" swimtime="00:01:26.97" resultid="4420" heatid="6152" lane="1" entrytime="00:01:26.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="233" reactiontime="+87" swimtime="00:03:19.70" resultid="4421" heatid="6270" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                    <SPLIT distance="100" swimtime="00:01:35.53" />
                    <SPLIT distance="150" swimtime="00:02:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="261" reactiontime="+88" swimtime="00:03:41.91" resultid="4422" heatid="6294" lane="3" entrytime="00:03:38.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.61" />
                    <SPLIT distance="100" swimtime="00:01:51.36" />
                    <SPLIT distance="150" swimtime="00:02:53.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="278" reactiontime="+111" swimtime="00:06:47.25" resultid="4423" heatid="6555" lane="5" entrytime="00:07:10.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.50" />
                    <SPLIT distance="100" swimtime="00:01:33.27" />
                    <SPLIT distance="150" swimtime="00:02:25.22" />
                    <SPLIT distance="200" swimtime="00:03:17.71" />
                    <SPLIT distance="250" swimtime="00:04:10.24" />
                    <SPLIT distance="300" swimtime="00:05:04.09" />
                    <SPLIT distance="350" swimtime="00:05:57.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-21" firstname="Marianna" gender="F" lastname="Michalczyk" nation="POL" athleteid="4424">
              <RESULTS>
                <RESULT eventid="1183" points="515" reactiontime="+83" swimtime="00:03:16.88" resultid="4425" heatid="6106" lane="6" entrytime="00:03:27.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                    <SPLIT distance="100" swimtime="00:01:35.14" />
                    <SPLIT distance="150" swimtime="00:02:26.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="480" reactiontime="+81" swimtime="00:01:13.34" resultid="4426" heatid="6155" lane="5" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="556" reactiontime="+87" swimtime="00:00:35.43" resultid="4427" heatid="6221" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1452" points="516" reactiontime="+75" swimtime="00:02:56.96" resultid="4428" heatid="6297" lane="6" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:25.70" />
                    <SPLIT distance="150" swimtime="00:02:17.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="4429" heatid="6337" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1595" points="468" reactiontime="+81" swimtime="00:01:31.02" resultid="4430" heatid="6508" lane="1" entrytime="00:01:35.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="4431">
              <RESULTS>
                <RESULT eventid="1228" points="683" reactiontime="+80" swimtime="00:00:29.68" resultid="4432" heatid="6138" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1272" points="697" reactiontime="+78" swimtime="00:00:57.03" resultid="4433" heatid="6179" lane="6" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="694" reactiontime="+80" swimtime="00:00:28.64" resultid="4434" heatid="6239" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="4435" heatid="6364" lane="1" entrytime="00:00:25.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="4436">
              <RESULTS>
                <RESULT eventid="1122" points="339" swimtime="00:17:13.76" resultid="4437" heatid="6442" lane="4" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.00" />
                    <SPLIT distance="100" swimtime="00:02:01.00" />
                    <SPLIT distance="150" swimtime="00:03:08.00" />
                    <SPLIT distance="200" swimtime="00:04:15.00" />
                    <SPLIT distance="250" swimtime="00:05:20.00" />
                    <SPLIT distance="300" swimtime="00:06:25.00" />
                    <SPLIT distance="350" swimtime="00:07:30.00" />
                    <SPLIT distance="400" swimtime="00:08:36.00" />
                    <SPLIT distance="450" swimtime="00:09:41.00" />
                    <SPLIT distance="500" swimtime="00:10:45.00" />
                    <SPLIT distance="550" swimtime="00:11:53.00" />
                    <SPLIT distance="600" swimtime="00:12:57.00" />
                    <SPLIT distance="650" swimtime="00:14:00.00" />
                    <SPLIT distance="700" swimtime="00:15:07.00" />
                    <SPLIT distance="750" swimtime="00:16:11.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="279" reactiontime="+102" swimtime="00:01:49.20" resultid="4438" heatid="6149" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="304" reactiontime="+83" swimtime="00:04:00.78" resultid="4439" heatid="6271" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.72" />
                    <SPLIT distance="100" swimtime="00:01:54.13" />
                    <SPLIT distance="150" swimtime="00:02:59.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="308" reactiontime="+97" swimtime="00:00:47.60" resultid="4440" heatid="6329" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1625" points="311" reactiontime="+106" swimtime="00:08:27.52" resultid="4441" heatid="6554" lane="4" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.17" />
                    <SPLIT distance="100" swimtime="00:02:00.27" />
                    <SPLIT distance="200" swimtime="00:04:13.21" />
                    <SPLIT distance="300" swimtime="00:06:25.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-04" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="4442">
              <RESULTS>
                <RESULT eventid="1168" points="854" reactiontime="+80" swimtime="00:01:01.40" resultid="4443" heatid="6100" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="828" reactiontime="+79" swimtime="00:00:26.89" resultid="4444" heatid="6240" lane="1" entrytime="00:00:27.80" />
                <RESULT comment="Rekord Polski kat. B" eventid="1528" points="858" reactiontime="+78" swimtime="00:00:24.27" resultid="4445" heatid="6365" lane="4" entrytime="00:00:24.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-13" firstname="Agnieszka" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="4446">
              <RESULTS>
                <RESULT eventid="1153" points="382" reactiontime="+85" swimtime="00:01:29.61" resultid="4447" heatid="6078" lane="5" entrytime="00:01:30.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="368" reactiontime="+84" swimtime="00:01:21.02" resultid="4448" heatid="6153" lane="4" entrytime="00:01:21.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="384" reactiontime="+106" swimtime="00:03:16.50" resultid="4449" heatid="6295" lane="4" entrytime="00:03:18.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                    <SPLIT distance="100" swimtime="00:01:34.89" />
                    <SPLIT distance="150" swimtime="00:02:30.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="348" reactiontime="+99" swimtime="00:06:20.99" resultid="4450" heatid="6555" lane="3" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                    <SPLIT distance="100" swimtime="00:01:31.12" />
                    <SPLIT distance="150" swimtime="00:02:19.26" />
                    <SPLIT distance="200" swimtime="00:03:08.10" />
                    <SPLIT distance="250" swimtime="00:03:57.31" />
                    <SPLIT distance="300" swimtime="00:04:46.60" />
                    <SPLIT distance="350" swimtime="00:05:35.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-12-31" firstname="Anna" gender="F" lastname="Michalska" nation="POL" athleteid="4451">
              <RESULTS>
                <RESULT eventid="1183" points="514" reactiontime="+113" swimtime="00:03:33.59" resultid="4452" heatid="6105" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.12" />
                    <SPLIT distance="100" swimtime="00:01:43.09" />
                    <SPLIT distance="150" swimtime="00:02:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="497" swimtime="00:00:45.54" resultid="4453" heatid="6198" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1422" points="266" swimtime="00:03:34.46" resultid="4454" heatid="6273" lane="2" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                    <SPLIT distance="100" swimtime="00:01:43.29" />
                    <SPLIT distance="150" swimtime="00:02:39.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="490" reactiontime="+93" swimtime="00:01:40.55" resultid="4455" heatid="6507" lane="5" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-03-16" firstname="Ewa" gender="F" lastname="Kosmol" nation="POL" athleteid="4456">
              <RESULTS>
                <RESULT eventid="1153" status="DNS" swimtime="00:00:00.00" resultid="4457" heatid="6076" lane="1" entrytime="00:01:45.00" />
                <RESULT eventid="1257" status="DNS" swimtime="00:00:00.00" resultid="4458" heatid="6150" lane="4" entrytime="00:01:40.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="4459" heatid="6272" lane="1" entrytime="00:03:45.00" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="4460" heatid="6332" lane="6" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisřaw" gender="M" lastname="Kozak" nation="POL" athleteid="4462">
              <RESULTS>
                <RESULT eventid="1198" points="643" reactiontime="+98" swimtime="00:02:44.41" resultid="4463" heatid="6117" lane="1" entrytime="00:02:39.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:18.78" />
                    <SPLIT distance="150" swimtime="00:02:02.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="720" swimtime="00:00:31.55" resultid="4464" heatid="6217" lane="2" entrytime="00:00:30.46" />
                <RESULT eventid="1363" points="595" reactiontime="+96" swimtime="00:00:30.15" resultid="4465" heatid="6236" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1610" points="739" reactiontime="+94" swimtime="00:01:09.89" resultid="4466" heatid="6408" lane="4" entrytime="00:01:07.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-22" firstname="Karol" gender="M" lastname="Dzięcioł" nation="POL" athleteid="4467">
              <RESULTS>
                <RESULT eventid="1272" points="743" reactiontime="+74" swimtime="00:00:55.91" resultid="4468" heatid="6179" lane="5" entrytime="00:00:56.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="614" reactiontime="+72" swimtime="00:00:27.14" resultid="4469" heatid="6364" lane="3" entrytime="00:00:25.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-17" firstname="Marek" gender="M" lastname="Makay" nation="POL" athleteid="4470">
              <RESULTS>
                <RESULT eventid="1137" points="668" swimtime="00:11:34.34" resultid="4471" heatid="6452" lane="2" entrytime="00:11:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:20.95" />
                    <SPLIT distance="200" swimtime="00:02:46.86" />
                    <SPLIT distance="300" swimtime="00:04:13.75" />
                    <SPLIT distance="400" swimtime="00:05:41.96" />
                    <SPLIT distance="500" swimtime="00:07:10.64" />
                    <SPLIT distance="600" swimtime="00:08:39.65" />
                    <SPLIT distance="700" swimtime="00:10:07.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="613" reactiontime="+71" swimtime="00:00:39.36" resultid="4472" heatid="6131" lane="5" entrytime="00:00:39.50" />
                <RESULT eventid="1272" points="732" swimtime="00:01:09.19" resultid="4473" heatid="6167" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="644" reactiontime="+77" swimtime="00:01:25.21" resultid="4474" heatid="6255" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="750" reactiontime="+115" swimtime="00:02:35.40" resultid="4475" heatid="6284" lane="1" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:01:14.45" />
                    <SPLIT distance="150" swimtime="00:01:55.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="648" reactiontime="+72" swimtime="00:03:07.02" resultid="4476" heatid="6376" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="100" swimtime="00:01:29.22" />
                    <SPLIT distance="150" swimtime="00:02:18.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="666" reactiontime="+113" swimtime="00:05:37.85" resultid="4477" heatid="6564" lane="3" entrytime="00:05:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:21.49" />
                    <SPLIT distance="150" swimtime="00:02:05.59" />
                    <SPLIT distance="200" swimtime="00:02:49.41" />
                    <SPLIT distance="250" swimtime="00:03:32.62" />
                    <SPLIT distance="300" swimtime="00:04:15.48" />
                    <SPLIT distance="350" swimtime="00:04:57.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-24" firstname="Ewa" gender="F" lastname="Szlagor" nation="POL" athleteid="4478">
              <RESULTS>
                <RESULT eventid="1153" points="768" reactiontime="+83" swimtime="00:01:14.64" resultid="4479" heatid="6082" lane="2" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="877" reactiontime="+78" swimtime="00:00:35.53" resultid="4480" heatid="6192" lane="5" />
                <RESULT eventid="1348" points="872" reactiontime="+82" swimtime="00:00:31.04" resultid="4481" heatid="6223" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1513" points="803" reactiontime="+81" swimtime="00:00:29.26" resultid="4482" heatid="6340" lane="5" entrytime="00:00:29.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1250" status="DNS" swimtime="00:00:00.00" resultid="4486" heatid="6525" lane="3" entrytime="00:02:01.12">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4330" number="1" />
                    <RELAYPOSITION athleteid="4304" number="2" />
                    <RELAYPOSITION athleteid="4392" number="3" />
                    <RELAYPOSITION athleteid="4359" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+85" swimtime="00:02:44.19" resultid="4487" heatid="6522" lane="5" entrytime="00:02:42.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                    <SPLIT distance="100" swimtime="00:01:33.92" />
                    <SPLIT distance="150" swimtime="00:02:14.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4322" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="4402" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4346" number="3" reactiontime="+8" />
                    <RELAYPOSITION athleteid="4352" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="6">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. B" eventid="1250" reactiontime="+65" swimtime="00:01:50.49" resultid="4488" heatid="6526" lane="4" entrytime="00:01:49.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.29" />
                    <SPLIT distance="100" swimtime="00:00:58.71" />
                    <SPLIT distance="150" swimtime="00:01:25.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4316" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="4462" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="4442" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4467" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+82" swimtime="00:01:41.62" resultid="4490" heatid="6534" lane="4" entrytime="00:01:44.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.76" />
                    <SPLIT distance="100" swimtime="00:00:52.92" />
                    <SPLIT distance="150" swimtime="00:01:17.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4311" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="4392" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4431" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="4442" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+94" swimtime="00:01:57.06" resultid="4491" heatid="6532" lane="3" entrytime="00:01:56.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                    <SPLIT distance="100" swimtime="00:00:58.08" />
                    <SPLIT distance="150" swimtime="00:01:27.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4330" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="4462" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="4352" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4359" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="10">
              <RESULTS>
                <RESULT eventid="1415" reactiontime="+96" swimtime="00:02:31.33" resultid="4492" heatid="6530" lane="3" entrytime="00:02:25.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="100" swimtime="00:01:16.82" />
                    <SPLIT distance="150" swimtime="00:01:54.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4365" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="4322" number="2" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4402" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4346" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1243" reactiontime="+73" swimtime="00:02:27.77" resultid="4485" heatid="6520" lane="5" entrytime="00:02:29.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="150" swimtime="00:01:49.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4410" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4478" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="4424" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4417" number="4" reactiontime="+98" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="7">
              <RESULTS>
                <RESULT eventid="1408" reactiontime="+54" swimtime="00:02:13.39" resultid="4489" heatid="6528" lane="2" entrytime="00:02:13.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:05.67" />
                    <SPLIT distance="150" swimtime="00:01:44.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4424" number="1" reactiontime="+54" />
                    <RELAYPOSITION athleteid="4410" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="4417" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="4478" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+81" swimtime="00:02:10.54" resultid="4483" heatid="6496" lane="2" entrytime="00:02:10.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:08.14" />
                    <SPLIT distance="150" swimtime="00:01:43.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4410" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4446" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="4346" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="4392" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1107" reactiontime="+96" swimtime="00:02:33.65" resultid="4484" heatid="6495" lane="5" entrytime="00:02:33.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="150" swimtime="00:01:59.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4417" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="4451" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="4322" number="3" />
                    <RELAYPOSITION athleteid="4402" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="11">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+82" swimtime="00:02:17.37" resultid="4493" heatid="6537" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                    <SPLIT distance="100" swimtime="00:01:14.87" />
                    <SPLIT distance="150" swimtime="00:01:44.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4442" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="4451" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4330" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="4410" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="12">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+82" swimtime="00:02:14.69" resultid="4494" heatid="6537" lane="3" entrytime="00:02:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                    <SPLIT distance="100" swimtime="00:01:11.85" />
                    <SPLIT distance="150" swimtime="00:01:42.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4431" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="4424" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="4392" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="4297" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="13">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+82" swimtime="00:02:44.02" resultid="4495" heatid="6536" lane="6" entrytime="00:02:45.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:25.60" />
                    <SPLIT distance="150" swimtime="00:02:05.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4352" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="4446" number="2" reactiontime="+84" />
                    <RELAYPOSITION athleteid="4346" number="3" reactiontime="+9" />
                    <RELAYPOSITION athleteid="4417" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Aquapark Wrocław" nation="POL" region="DOL">
          <CONTACT city="Wrocław" name="Stasiaczek" phone="792883772" street="Sztabowa 78/10" zip="53-310" />
          <ATHLETES>
            <ATHLETE birthdate="1990-04-04" firstname="Krystian" gender="M" lastname="Lipowczyk" nation="POL" athleteid="4528">
              <RESULTS>
                <RESULT eventid="1168" points="561" reactiontime="+71" swimtime="00:01:11.75" resultid="4529" heatid="6093" lane="4" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="524" reactiontime="+73" swimtime="00:01:01.22" resultid="4530" heatid="6170" lane="6" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="363" reactiontime="+76" swimtime="00:01:16.20" resultid="4531" heatid="6260" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="4532" heatid="6357" lane="1" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-21" firstname="Mateusz" gender="M" lastname="Dudek" nation="POL" athleteid="4533">
              <RESULTS>
                <RESULT eventid="1198" points="668" reactiontime="+77" swimtime="00:02:34.19" resultid="4534" heatid="6117" lane="4" entrytime="00:02:32.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:12.88" />
                    <SPLIT distance="150" swimtime="00:01:53.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="748" reactiontime="+74" swimtime="00:00:31.20" resultid="4535" heatid="6216" lane="3" entrytime="00:00:31.80" />
                <RESULT eventid="1610" points="705" reactiontime="+74" swimtime="00:01:09.83" resultid="4536" heatid="6408" lane="5" entrytime="00:01:09.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-09" firstname="Paweł" gender="M" lastname="Handke" nation="POL" athleteid="4537">
              <RESULTS>
                <RESULT eventid="1198" points="649" reactiontime="+84" swimtime="00:02:43.92" resultid="4538" heatid="6117" lane="5" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:19.16" />
                    <SPLIT distance="150" swimtime="00:02:01.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="743" reactiontime="+78" swimtime="00:00:55.83" resultid="4539" heatid="6179" lane="3" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="4540" heatid="6292" lane="5" entrytime="00:02:04.00" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="4541" heatid="6365" lane="3" entrytime="00:00:24.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-04-29" firstname="Łukasz" gender="M" lastname="Lesiewicz" nation="POL" athleteid="4543">
              <RESULTS>
                <RESULT eventid="1168" reactiontime="+82" status="DNF" swimtime="00:00:00.00" resultid="4544" heatid="6097" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="543" reactiontime="+66" swimtime="00:00:31.19" resultid="4545" heatid="6138" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1393" points="504" reactiontime="+67" swimtime="00:01:08.30" resultid="4546" heatid="6261" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="4547" heatid="6363" lane="5" entrytime="00:00:26.00" />
                <RESULT eventid="1558" points="480" reactiontime="+61" swimtime="00:02:35.41" resultid="4548" heatid="6380" lane="5" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                    <SPLIT distance="150" swimtime="00:01:55.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-10" firstname="Jarosław" gender="M" lastname="Wnęk" nation="POL" athleteid="4549">
              <RESULTS>
                <RESULT eventid="1137" points="404" swimtime="00:11:10.82" resultid="4550" heatid="6457" lane="2" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:08.40" />
                    <SPLIT distance="200" swimtime="00:02:25.04" />
                    <SPLIT distance="300" swimtime="00:03:46.03" />
                    <SPLIT distance="400" swimtime="00:05:09.54" />
                    <SPLIT distance="500" swimtime="00:06:39.74" />
                    <SPLIT distance="600" swimtime="00:08:09.95" />
                    <SPLIT distance="700" swimtime="00:09:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="324" reactiontime="+88" swimtime="00:02:54.71" resultid="4551" heatid="6188" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:17.94" />
                    <SPLIT distance="150" swimtime="00:02:03.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" status="DNS" swimtime="00:00:00.00" resultid="4552" heatid="6569" lane="2" entrytime="00:04:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-11-17" firstname="Michał" gender="M" lastname="Stasiaczek" nation="POL" athleteid="4553">
              <RESULTS>
                <RESULT eventid="1168" points="770" reactiontime="+80" swimtime="00:01:03.17" resultid="4554" heatid="6100" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="791" reactiontime="+76" swimtime="00:02:33.50" resultid="4555" heatid="6117" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:14.89" />
                    <SPLIT distance="150" swimtime="00:01:54.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="727" reactiontime="+76" swimtime="00:00:31.46" resultid="4556" heatid="6217" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="4557" heatid="6311" lane="2" entrytime="00:02:19.00" />
                <RESULT eventid="1610" points="798" reactiontime="+80" swimtime="00:01:08.11" resultid="4558" heatid="6408" lane="2" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" name="AZS AWF Katowice" nation="POL" region="SLA">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501 370 222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1991-09-13" firstname="Tomasz" gender="M" lastname="Czermak" nation="POL" license="S00611200197" athleteid="4560">
              <RESULTS>
                <RESULT eventid="1137" points="664" swimtime="00:09:28.62" resultid="4561" heatid="6457" lane="4" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:05.62" />
                    <SPLIT distance="200" swimtime="00:02:14.74" />
                    <SPLIT distance="300" swimtime="00:03:25.76" />
                    <SPLIT distance="400" swimtime="00:04:37.53" />
                    <SPLIT distance="500" swimtime="00:05:50.29" />
                    <SPLIT distance="600" swimtime="00:07:03.87" />
                    <SPLIT distance="700" swimtime="00:08:17.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="707" reactiontime="+75" swimtime="00:02:31.37" resultid="4562" heatid="6117" lane="3" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:12.71" />
                    <SPLIT distance="150" swimtime="00:01:52.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="527" reactiontime="+74" swimtime="00:02:28.54" resultid="4563" heatid="6191" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:10.72" />
                    <SPLIT distance="150" swimtime="00:01:49.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="748" reactiontime="+72" swimtime="00:00:31.20" resultid="4564" heatid="6217" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1467" points="656" reactiontime="+74" swimtime="00:02:22.04" resultid="4565" heatid="6311" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:10.05" />
                    <SPLIT distance="150" swimtime="00:01:49.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="712" reactiontime="+73" swimtime="00:01:09.60" resultid="4566" heatid="6408" lane="3" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="626" reactiontime="+71" swimtime="00:04:32.27" resultid="4567" heatid="6570" lane="5" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:04.12" />
                    <SPLIT distance="150" swimtime="00:01:38.50" />
                    <SPLIT distance="200" swimtime="00:02:13.19" />
                    <SPLIT distance="250" swimtime="00:02:48.37" />
                    <SPLIT distance="300" swimtime="00:03:23.43" />
                    <SPLIT distance="350" swimtime="00:03:58.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-10-04" firstname="Kuba" gender="M" lastname="Kowalik" nation="POL" athleteid="4618">
              <RESULTS>
                <RESULT eventid="1272" points="605" reactiontime="+72" swimtime="00:00:58.36" resultid="4619" heatid="6176" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="599" swimtime="00:00:29.43" resultid="4620" heatid="6238" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1437" points="446" reactiontime="+78" swimtime="00:02:20.87" resultid="4621" heatid="6287" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:04.68" />
                    <SPLIT distance="150" swimtime="00:01:42.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="584" reactiontime="+75" swimtime="00:00:26.70" resultid="4622" heatid="6360" lane="6" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UCWAR" name="UCSiR Warszawa" nation="POL" region="WAR">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1985-05-26" firstname="URSZULA" gender="F" lastname="BIELAWSKA" nation="POL" athleteid="4569">
              <RESULTS>
                <RESULT eventid="1122" points="438" swimtime="00:12:11.40" resultid="4570" heatid="6444" lane="5" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.44" />
                    <SPLIT distance="200" swimtime="00:02:53.48" />
                    <SPLIT distance="300" swimtime="00:04:27.91" />
                    <SPLIT distance="400" swimtime="00:06:01.55" />
                    <SPLIT distance="500" swimtime="00:07:35.75" />
                    <SPLIT distance="600" swimtime="00:09:09.32" />
                    <SPLIT distance="700" swimtime="00:10:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="406" reactiontime="+87" swimtime="00:01:28.56" resultid="4571" heatid="6079" lane="4" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="524" reactiontime="+83" swimtime="00:01:11.25" resultid="4572" heatid="6156" lane="3" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="487" reactiontime="+84" swimtime="00:00:43.31" resultid="4573" heatid="6199" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1422" points="456" reactiontime="+89" swimtime="00:02:39.62" resultid="4574" heatid="6276" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                    <SPLIT distance="150" swimtime="00:01:57.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="400" reactiontime="+76" swimtime="00:01:35.96" resultid="4575" heatid="6509" lane="6" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="461" reactiontime="+84" swimtime="00:05:44.23" resultid="4576" heatid="6557" lane="4" entrytime="00:05:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:20.41" />
                    <SPLIT distance="150" swimtime="00:02:03.95" />
                    <SPLIT distance="200" swimtime="00:02:48.29" />
                    <SPLIT distance="250" swimtime="00:03:32.85" />
                    <SPLIT distance="300" swimtime="00:04:17.97" />
                    <SPLIT distance="350" swimtime="00:05:02.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-05-26" firstname="MAŁGORZATA" gender="F" lastname="KOTAŃSKA" nation="POL" athleteid="4577">
              <RESULTS>
                <RESULT eventid="1122" points="336" swimtime="00:14:46.31" resultid="4578" heatid="6443" lane="1" entrytime="00:14:45.00" />
                <RESULT eventid="1183" points="536" reactiontime="+88" swimtime="00:03:30.63" resultid="4579" heatid="6105" lane="2" entrytime="00:03:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.60" />
                    <SPLIT distance="100" swimtime="00:01:40.34" />
                    <SPLIT distance="150" swimtime="00:02:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="423" reactiontime="+87" swimtime="00:01:24.58" resultid="4580" heatid="6153" lane="5" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="579" reactiontime="+97" swimtime="00:00:43.27" resultid="4581" heatid="6198" lane="3" entrytime="00:00:44.00" />
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="4582" heatid="6273" lane="3" entrytime="00:03:25.00" />
                <RESULT eventid="1513" points="407" reactiontime="+94" swimtime="00:00:37.98" resultid="4583" heatid="6333" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1595" points="595" reactiontime="+88" swimtime="00:01:34.22" resultid="4584" heatid="6508" lane="6" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="MICHAŁ" gender="M" lastname="NOWAK" nation="POL" athleteid="4585">
              <RESULTS>
                <RESULT eventid="1092" points="680" reactiontime="+94" swimtime="00:06:35.86" resultid="4586" heatid="6488" lane="5" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:01:34.80" />
                    <SPLIT distance="200" swimtime="00:03:19.57" />
                    <SPLIT distance="250" swimtime="00:04:11.97" />
                    <SPLIT distance="300" swimtime="00:05:02.95" />
                    <SPLIT distance="350" swimtime="00:05:50.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="774" reactiontime="+89" swimtime="00:01:18.29" resultid="4587" heatid="6090" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="880" reactiontime="+93" swimtime="00:03:04.20" resultid="4588" heatid="6113" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                    <SPLIT distance="100" swimtime="00:01:30.16" />
                    <SPLIT distance="150" swimtime="00:02:18.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="849" reactiontime="+94" swimtime="00:00:36.17" resultid="4589" heatid="6212" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1467" points="717" reactiontime="+95" swimtime="00:02:59.96" resultid="4590" heatid="6304" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:31.99" />
                    <SPLIT distance="150" swimtime="00:02:19.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="4591" heatid="6319" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1610" points="889" reactiontime="+90" swimtime="00:01:22.13" resultid="4592" heatid="6403" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CZEST" name="Częstochowa" nation="POL" region="SLA">
          <CONTACT name="Krogulec" />
          <ATHLETES>
            <ATHLETE birthdate="1981-11-02" firstname="Monika" gender="F" lastname="Nowak" nation="POL" athleteid="4596">
              <RESULTS>
                <RESULT eventid="1153" points="505" reactiontime="+91" swimtime="00:01:21.62" resultid="4597" heatid="6081" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="604" reactiontime="+89" swimtime="00:01:08.67" resultid="4598" heatid="6157" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="474" reactiontime="+91" swimtime="00:00:42.66" resultid="4599" heatid="6200" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="1422" points="533" reactiontime="+88" swimtime="00:02:34.45" resultid="4600" heatid="6276" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:01:54.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" reactiontime="+87" status="DNS" swimtime="00:00:00.00" resultid="4601" heatid="6339" lane="1" entrytime="00:00:30.50" />
                <RESULT eventid="1543" points="464" reactiontime="+81" swimtime="00:02:59.58" resultid="4602" heatid="6370" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:27.66" />
                    <SPLIT distance="150" swimtime="00:02:13.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-26" firstname="Rafał" gender="M" lastname="Nowak" nation="POL" athleteid="4603">
              <RESULTS>
                <RESULT eventid="1168" points="279" reactiontime="+87" swimtime="00:01:29.31" resultid="4604" heatid="6086" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="304" reactiontime="+86" swimtime="00:01:16.42" resultid="4605" heatid="6163" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="270" reactiontime="+98" swimtime="00:00:38.88" resultid="4606" heatid="6229" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1467" points="263" reactiontime="+89" swimtime="00:03:15.58" resultid="4607" heatid="6303" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                    <SPLIT distance="100" swimtime="00:01:32.60" />
                    <SPLIT distance="150" swimtime="00:02:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="4608" heatid="6319" lane="6" entrytime="00:01:30.00" />
                <RESULT eventid="1528" points="301" reactiontime="+88" swimtime="00:00:34.53" resultid="4609" heatid="6349" lane="4" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-07-31" firstname="Piotr" gender="M" lastname="Krogulec" nation="POL" athleteid="4610">
              <RESULTS>
                <RESULT eventid="1092" points="493" reactiontime="+85" swimtime="00:05:34.19" resultid="4611" heatid="6490" lane="6" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                    <SPLIT distance="100" swimtime="00:01:08.44" />
                    <SPLIT distance="150" swimtime="00:01:48.90" />
                    <SPLIT distance="200" swimtime="00:02:31.71" />
                    <SPLIT distance="250" swimtime="00:03:18.89" />
                    <SPLIT distance="300" swimtime="00:04:09.35" />
                    <SPLIT distance="350" swimtime="00:04:52.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="735" reactiontime="+81" swimtime="00:01:05.58" resultid="4612" heatid="6095" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="587" reactiontime="+63" swimtime="00:00:30.39" resultid="4613" heatid="6134" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1393" points="541" reactiontime="+72" swimtime="00:01:06.71" resultid="4614" heatid="6258" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="594" reactiontime="+78" swimtime="00:02:26.85" resultid="4615" heatid="6307" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:51.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="619" reactiontime="+74" swimtime="00:01:02.94" resultid="4616" heatid="6324" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="590" reactiontime="+73" swimtime="00:02:25.14" resultid="4617" heatid="6379" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:49.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="UKS Wodnik 29 Katowice" nation="POL">
          <CONTACT city="Katowice" email="bozenakaspmroz@o2.pl" name="Bożena Mrozińska" phone="502 013 302" street="Barbary 14/9" zip="40-053" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="4624">
              <RESULTS>
                <RESULT eventid="1198" points="646" reactiontime="+89" swimtime="00:03:06.47" resultid="4625" heatid="6113" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:01:30.36" />
                    <SPLIT distance="150" swimtime="00:02:18.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="4626" heatid="6175" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="754" reactiontime="+83" swimtime="00:00:35.37" resultid="4627" heatid="6213" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="4628" heatid="6305" lane="6" entrytime="00:02:55.00" />
                <RESULT eventid="1528" points="514" reactiontime="+82" swimtime="00:00:31.67" resultid="4629" heatid="6350" lane="3" entrytime="00:00:31.00" />
                <RESULT comment="K13" eventid="1610" reactiontime="+85" status="DSQ" swimtime="00:01:21.06" resultid="4630" heatid="6404" lane="4" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-05" firstname="Marcin" gender="M" lastname="Szczypiński" nation="POL" athleteid="4631">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. A" eventid="1137" points="779" swimtime="00:09:07.72" resultid="4632" heatid="6457" lane="5" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.08" />
                    <SPLIT distance="200" swimtime="00:02:11.50" />
                    <SPLIT distance="300" swimtime="00:03:21.15" />
                    <SPLIT distance="400" swimtime="00:04:30.56" />
                    <SPLIT distance="500" swimtime="00:05:39.50" />
                    <SPLIT distance="600" swimtime="00:06:48.19" />
                    <SPLIT distance="700" swimtime="00:07:58.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="804" reactiontime="+80" swimtime="00:00:54.39" resultid="4633" heatid="6180" lane="2" entrytime="00:00:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="750" reactiontime="+90" swimtime="00:02:18.52" resultid="4634" heatid="6191" lane="3" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:07.22" />
                    <SPLIT distance="150" swimtime="00:01:43.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="854" reactiontime="+57" swimtime="00:00:26.72" resultid="4635" heatid="6241" lane="2" entrytime="00:00:26.50" />
                <RESULT eventid="1437" points="765" reactiontime="+82" swimtime="00:02:01.01" resultid="4636" heatid="6292" lane="2" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="100" swimtime="00:00:58.21" />
                    <SPLIT distance="150" swimtime="00:01:29.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="836" reactiontime="+79" swimtime="00:00:58.96" resultid="4637" heatid="6327" lane="1" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" points="765" reactiontime="+80" swimtime="00:04:23.90" resultid="4638" heatid="6570" lane="2" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="100" swimtime="00:01:01.77" />
                    <SPLIT distance="150" swimtime="00:01:35.42" />
                    <SPLIT distance="200" swimtime="00:02:09.79" />
                    <SPLIT distance="250" swimtime="00:02:43.93" />
                    <SPLIT distance="300" swimtime="00:03:17.87" />
                    <SPLIT distance="350" swimtime="00:03:51.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-09" firstname="Krystyna" gender="F" lastname="Nicpoń" nation="POL" athleteid="4639">
              <RESULTS>
                <RESULT eventid="1153" points="404" reactiontime="+101" swimtime="00:02:10.69" resultid="4640" heatid="6075" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="525" reactiontime="+85" swimtime="00:00:53.96" resultid="4641" heatid="6120" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="1378" points="670" reactiontime="+77" swimtime="00:01:55.65" resultid="4642" heatid="6244" lane="3" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="685" reactiontime="+79" swimtime="00:04:08.15" resultid="4643" heatid="6367" lane="3" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.89" />
                    <SPLIT distance="100" swimtime="00:01:56.66" />
                    <SPLIT distance="150" swimtime="00:03:02.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-05-18" firstname="Urszula" gender="F" lastname="Walkowicz" nation="POL" athleteid="4644">
              <RESULTS>
                <RESULT eventid="1122" points="328" swimtime="00:24:53.86" resultid="4645" heatid="6441" lane="4" entrytime="00:22:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.95" />
                    <SPLIT distance="150" swimtime="00:02:44.86" />
                    <SPLIT distance="250" swimtime="00:05:45.89" />
                    <SPLIT distance="300" swimtime="00:08:54.67" />
                    <SPLIT distance="400" swimtime="00:12:07.16" />
                    <SPLIT distance="500" swimtime="00:15:19.95" />
                    <SPLIT distance="600" swimtime="00:18:34.36" />
                    <SPLIT distance="700" swimtime="00:21:54.64" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski kat. L" eventid="1213" points="503" reactiontime="+77" swimtime="00:01:09.27" resultid="4646" heatid="6119" lane="2" entrytime="00:01:05.00" />
                <RESULT comment="Rekord Polski kat. L" eventid="1378" points="576" reactiontime="+79" swimtime="00:02:36.91" resultid="4647" heatid="6243" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="363" reactiontime="+106" swimtime="00:01:03.04" resultid="4648" heatid="6329" lane="4" entrytime="00:01:05.00" />
                <RESULT comment="Rekord Polski kat. L" eventid="1543" points="570" reactiontime="+71" swimtime="00:05:45.33" resultid="4649" heatid="6367" lane="5" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.37" />
                    <SPLIT distance="100" swimtime="00:02:51.85" />
                    <SPLIT distance="150" swimtime="00:04:21.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-02-02" firstname="Maria" gender="F" lastname="Śmiglewska" nation="POL" athleteid="4650">
              <RESULTS>
                <RESULT eventid="1183" points="209" swimtime="00:07:08.86" resultid="4651" heatid="6101" lane="3" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:43.36" />
                    <SPLIT distance="100" swimtime="00:03:30.52" />
                    <SPLIT distance="150" swimtime="00:05:23.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="268" reactiontime="+138" swimtime="00:01:14.36" resultid="4652" heatid="6118" lane="2" entrytime="00:01:25.00" />
                <RESULT eventid="1318" points="119" swimtime="00:01:35.61" resultid="4653" heatid="6192" lane="3" entrytime="00:01:35.00" />
                <RESULT eventid="1378" points="223" reactiontime="+130" swimtime="00:02:56.76" resultid="4654" heatid="6242" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="4655">
              <RESULTS>
                <RESULT eventid="1137" points="609" swimtime="00:10:49.07" resultid="4656" heatid="6454" lane="2" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:15.44" />
                    <SPLIT distance="200" swimtime="00:02:35.29" />
                    <SPLIT distance="300" swimtime="00:03:57.08" />
                    <SPLIT distance="400" swimtime="00:05:18.72" />
                    <SPLIT distance="500" swimtime="00:06:40.69" />
                    <SPLIT distance="600" swimtime="00:08:03.96" />
                    <SPLIT distance="700" swimtime="00:09:27.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="609" reactiontime="+74" swimtime="00:00:34.04" resultid="4657" heatid="6134" lane="6" entrytime="00:00:34.60" />
                <RESULT eventid="1272" points="663" reactiontime="+92" swimtime="00:01:02.79" resultid="4658" heatid="6171" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="701" reactiontime="+83" swimtime="00:01:13.24" resultid="4659" heatid="6257" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="671" reactiontime="+91" swimtime="00:02:20.00" resultid="4660" heatid="6287" lane="5" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                    <SPLIT distance="100" swimtime="00:01:07.42" />
                    <SPLIT distance="150" swimtime="00:01:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="681" reactiontime="+86" swimtime="00:00:27.88" resultid="4661" heatid="6354" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1558" points="701" reactiontime="+79" swimtime="00:02:38.61" resultid="4662" heatid="6377" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:17.76" />
                    <SPLIT distance="150" swimtime="00:01:58.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-04-23" firstname="Agata" gender="F" lastname="Wolińska" nation="POL" athleteid="4663">
              <RESULTS>
                <RESULT eventid="1153" points="187" reactiontime="+90" swimtime="00:02:05.22" resultid="4664" heatid="6075" lane="1" entrytime="00:02:02.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="187" reactiontime="+85" swimtime="00:01:50.90" resultid="4665" heatid="6149" lane="3" entrytime="00:01:48.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" points="109" reactiontime="+84" swimtime="00:01:03.73" resultid="4666" heatid="6218" lane="4" entrytime="00:00:58.61" />
                <RESULT eventid="1422" points="161" swimtime="00:04:13.29" resultid="4667" heatid="6270" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.12" />
                    <SPLIT distance="100" swimtime="00:01:53.21" />
                    <SPLIT distance="150" swimtime="00:03:02.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="220" reactiontime="+91" swimtime="00:00:46.60" resultid="4668" heatid="6331" lane="6" entrytime="00:00:44.64" />
                <RESULT eventid="1595" points="163" reactiontime="+98" swimtime="00:02:24.89" resultid="4669" heatid="6502" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-19" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="4670">
              <RESULTS>
                <RESULT eventid="1272" points="615" reactiontime="+87" swimtime="00:01:13.32" resultid="4671" heatid="6163" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="427" reactiontime="+92" swimtime="00:03:35.16" resultid="4672" heatid="6186" lane="6" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                    <SPLIT distance="100" swimtime="00:01:38.69" />
                    <SPLIT distance="150" swimtime="00:02:37.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-4 - przedwczesny start." eventid="1363" reactiontime="+74" status="DSQ" swimtime="00:00:34.12" resultid="4673" heatid="6230" lane="1" entrytime="00:00:33.50" />
                <RESULT eventid="1437" points="499" reactiontime="+98" swimtime="00:02:58.01" resultid="4674" heatid="6280" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                    <SPLIT distance="100" swimtime="00:01:25.29" />
                    <SPLIT distance="150" swimtime="00:02:14.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="563" reactiontime="+93" swimtime="00:01:24.82" resultid="4675" heatid="6320" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="587" reactiontime="+99" swimtime="00:00:32.58" resultid="4676" heatid="6348" lane="1" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-03-15" firstname="Jolanta" gender="F" lastname="Stefanek" nation="POL" athleteid="4677">
              <RESULTS>
                <RESULT eventid="1183" points="621" reactiontime="+81" swimtime="00:03:29.11" resultid="4678" heatid="6106" lane="1" entrytime="00:03:26.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.23" />
                    <SPLIT distance="100" swimtime="00:01:40.77" />
                    <SPLIT distance="150" swimtime="00:02:35.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="636" reactiontime="+81" swimtime="00:00:44.07" resultid="4679" heatid="6199" lane="1" entrytime="00:00:42.43" />
                <RESULT eventid="1452" points="395" reactiontime="+87" swimtime="00:03:42.25" resultid="4680" heatid="6295" lane="1" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.59" />
                    <SPLIT distance="100" swimtime="00:01:46.89" />
                    <SPLIT distance="150" swimtime="00:02:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="618" reactiontime="+84" swimtime="00:01:37.83" resultid="4681" heatid="6508" lane="2" entrytime="00:01:34.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="4682">
              <RESULTS>
                <RESULT eventid="1153" points="619" reactiontime="+88" swimtime="00:01:16.27" resultid="4683" heatid="6081" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="685" reactiontime="+80" swimtime="00:01:05.86" resultid="4684" heatid="6158" lane="6" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1348" status="DNS" swimtime="00:00:00.00" resultid="4685" heatid="6223" lane="5" entrytime="00:00:31.50" />
                <RESULT eventid="1452" status="DNS" swimtime="00:00:00.00" resultid="4686" heatid="6297" lane="3" entrytime="00:02:50.00" />
                <RESULT eventid="1483" status="DNS" swimtime="00:00:00.00" resultid="4687" heatid="6315" lane="5" entrytime="00:01:16.50" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="4688" heatid="6340" lane="1" entrytime="00:00:29.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-12-22" firstname="Sylwia" gender="F" lastname="Kornaś" nation="POL" athleteid="4689">
              <RESULTS>
                <RESULT eventid="1213" points="365" reactiontime="+76" swimtime="00:00:42.59" resultid="4690" heatid="6122" lane="2" entrytime="00:00:43.02" />
                <RESULT eventid="1257" points="364" reactiontime="+82" swimtime="00:01:20.41" resultid="4691" heatid="6152" lane="5" entrytime="00:01:26.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="399" reactiontime="+87" swimtime="00:00:46.29" resultid="4692" heatid="6197" lane="4" entrytime="00:00:47.66" />
                <RESULT eventid="1378" points="309" reactiontime="+72" swimtime="00:01:33.80" resultid="4693" heatid="6245" lane="4" entrytime="00:01:35.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="383" reactiontime="+80" swimtime="00:00:36.33" resultid="4694" heatid="6334" lane="2" entrytime="00:00:36.48" />
                <RESULT eventid="1543" points="309" reactiontime="+75" swimtime="00:03:19.90" resultid="4695" heatid="6368" lane="3" entrytime="00:03:25.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                    <SPLIT distance="100" swimtime="00:01:37.00" />
                    <SPLIT distance="150" swimtime="00:02:28.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-05-05" firstname="Marek" gender="M" lastname="Mróz" nation="POL" athleteid="4696">
              <RESULTS>
                <RESULT eventid="1137" points="581" swimtime="00:10:03.78" resultid="6500" heatid="6446" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:07.86" />
                    <SPLIT distance="200" swimtime="00:02:20.15" />
                    <SPLIT distance="300" swimtime="00:03:34.18" />
                    <SPLIT distance="400" swimtime="00:04:51.87" />
                    <SPLIT distance="500" swimtime="00:06:11.22" />
                    <SPLIT distance="600" swimtime="00:07:26.52" />
                    <SPLIT distance="700" swimtime="00:08:46.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="4698" heatid="6179" lane="2" entrytime="00:00:56.50" />
                <RESULT eventid="1363" points="790" reactiontime="+79" swimtime="00:00:27.43" resultid="4699" heatid="6240" lane="2" entrytime="00:00:27.30" />
                <RESULT eventid="1437" status="DNS" swimtime="00:00:00.00" resultid="4700" heatid="6290" lane="3" entrytime="00:02:10.00" />
                <RESULT eventid="1528" points="695" reactiontime="+78" swimtime="00:00:25.67" resultid="4701" heatid="6365" lane="6" entrytime="00:00:25.13" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-03-30" firstname="Mateusz" gender="M" lastname="Gawełczyk" nation="POL" athleteid="4702">
              <RESULTS>
                <RESULT eventid="1137" points="751" swimtime="00:09:05.62" resultid="4703" heatid="6457" lane="3" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:03.68" />
                    <SPLIT distance="200" swimtime="00:02:10.50" />
                    <SPLIT distance="300" swimtime="00:03:18.74" />
                    <SPLIT distance="400" swimtime="00:04:27.87" />
                    <SPLIT distance="500" swimtime="00:05:37.28" />
                    <SPLIT distance="600" swimtime="00:06:46.94" />
                    <SPLIT distance="700" swimtime="00:07:56.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" status="DNS" swimtime="00:00:00.00" resultid="4704" heatid="6570" lane="4" entrytime="00:04:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-16" firstname="Michał" gender="M" lastname="SPŁAWIŃSKI" nation="POL" athleteid="4705">
              <RESULTS>
                <RESULT eventid="1610" points="659" reactiontime="+81" swimtime="00:01:14.52" resultid="6571" heatid="6408" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="489" reactiontime="+94" swimtime="00:05:48.65" resultid="4706" heatid="6488" lane="6" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:18.92" />
                    <SPLIT distance="150" swimtime="00:02:04.63" />
                    <SPLIT distance="200" swimtime="00:02:52.11" />
                    <SPLIT distance="250" swimtime="00:03:39.92" />
                    <SPLIT distance="300" swimtime="00:04:25.56" />
                    <SPLIT distance="350" swimtime="00:05:08.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="659" reactiontime="+100" swimtime="00:01:06.96" resultid="4707" heatid="6094" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="594" reactiontime="+64" swimtime="00:00:31.05" resultid="4708" heatid="6137" lane="2" entrytime="00:00:30.50" />
                <RESULT eventid="1333" points="894" reactiontime="+78" swimtime="00:00:30.58" resultid="4709" heatid="6217" lane="1" entrytime="00:00:30.70" />
                <RESULT eventid="1363" points="808" reactiontime="+81" swimtime="00:00:27.12" resultid="4710" heatid="6241" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1528" points="789" reactiontime="+75" swimtime="00:00:24.96" resultid="4711" heatid="6365" lane="1" entrytime="00:00:25.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-05-08" firstname="Bartłomiej" gender="M" lastname="Kułaga" nation="POL" athleteid="4712">
              <RESULTS>
                <RESULT eventid="1302" points="598" reactiontime="+91" swimtime="00:02:29.31" resultid="4713" heatid="6190" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:08.81" />
                    <SPLIT distance="150" swimtime="00:01:47.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="683" reactiontime="+83" swimtime="00:00:28.68" resultid="4714" heatid="6240" lane="6" entrytime="00:00:27.80" />
                <RESULT eventid="1498" points="610" reactiontime="+82" swimtime="00:01:05.68" resultid="4715" heatid="6326" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="4716">
              <RESULTS>
                <RESULT eventid="1272" points="571" reactiontime="+93" swimtime="00:01:08.57" resultid="4717" heatid="6169" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="673" reactiontime="+91" swimtime="00:00:31.63" resultid="4718" heatid="6232" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1528" points="640" reactiontime="+93" swimtime="00:00:29.43" resultid="4719" heatid="6353" lane="3" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-11-14" firstname="Aleksander" gender="M" lastname="Aleksandrowicz" nation="POL" athleteid="4720">
              <RESULTS>
                <RESULT eventid="1228" points="333" reactiontime="+172" swimtime="00:00:57.00" resultid="4721" heatid="6129" lane="4" entrytime="00:00:45.00" />
                <RESULT comment="O-4" eventid="1333" status="DSQ" swimtime="00:01:01.17" resultid="4722" heatid="6203" lane="2" entrytime="00:00:55.00" />
                <RESULT eventid="1393" points="380" reactiontime="+93" swimtime="00:02:01.55" resultid="4723" heatid="6252" lane="6" entrytime="00:01:50.00" />
                <RESULT eventid="1528" points="504" reactiontime="+99" swimtime="00:00:41.18" resultid="4724" heatid="6343" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1610" points="292" reactiontime="+106" swimtime="00:02:13.52" resultid="4725" heatid="6395" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Olga" gender="F" lastname="Załuska" nation="POL" athleteid="4726">
              <RESULTS>
                <RESULT eventid="1348" points="544" reactiontime="+84" swimtime="00:00:33.79" resultid="4737" heatid="6223" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="4738" heatid="6338" lane="2" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski kat. B" eventid="1415" reactiontime="+79" swimtime="00:01:41.02" resultid="4729" heatid="6534" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.62" />
                    <SPLIT distance="100" swimtime="00:00:51.83" />
                    <SPLIT distance="150" swimtime="00:01:16.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4705" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4712" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4696" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="4631" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1250" reactiontime="+74" swimtime="00:01:52.19" resultid="4730" heatid="6526" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                    <SPLIT distance="100" swimtime="00:00:58.80" />
                    <SPLIT distance="150" swimtime="00:01:27.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4631" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4705" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="4712" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="4696" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1250" reactiontime="+81" swimtime="00:02:12.81" resultid="4735" heatid="6524" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:43.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4655" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4624" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4670" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="4716" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1415" reactiontime="+86" swimtime="00:02:00.37" resultid="4736" heatid="6532" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                    <SPLIT distance="100" swimtime="00:00:59.45" />
                    <SPLIT distance="150" swimtime="00:01:31.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4655" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="4624" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4670" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="4716" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1408" reactiontime="+86" swimtime="00:02:54.25" resultid="4731" heatid="6527" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.67" />
                    <SPLIT distance="100" swimtime="00:01:35.72" />
                    <SPLIT distance="150" swimtime="00:02:16.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4663" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="4639" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4677" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="4689" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1243" status="DNS" swimtime="00:00:00.00" resultid="4732" heatid="6519" lane="5" entrytime="00:03:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4639" number="1" />
                    <RELAYPOSITION athleteid="4677" number="2" />
                    <RELAYPOSITION athleteid="4682" number="3" />
                    <RELAYPOSITION athleteid="4689" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+76" swimtime="00:02:30.01" resultid="4733" heatid="6538" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                    <SPLIT distance="100" swimtime="00:01:15.80" />
                    <SPLIT distance="150" swimtime="00:01:43.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4689" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4705" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="4696" number="3" reactiontime="+8" />
                    <RELAYPOSITION athleteid="4663" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1588" reactiontime="+78" swimtime="00:02:42.91" resultid="4734" heatid="6536" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.96" />
                    <SPLIT distance="100" swimtime="00:01:37.62" />
                    <SPLIT distance="150" swimtime="00:02:12.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4639" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4677" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4670" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="4716" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01511" name="MTP Delfin Cieszyn" nation="POL" region="11">
          <ATHLETES>
            <ATHLETE birthdate="1990-06-12" firstname="Katarzyna" gender="F" lastname="Widzik" nation="POL" athleteid="4760">
              <RESULTS>
                <RESULT eventid="1058" points="432" reactiontime="+81" swimtime="00:06:24.21" resultid="4761" heatid="6428" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:01:31.70" />
                    <SPLIT distance="150" swimtime="00:02:18.91" />
                    <SPLIT distance="200" swimtime="00:03:05.22" />
                    <SPLIT distance="250" swimtime="00:04:00.14" />
                    <SPLIT distance="300" swimtime="00:04:55.25" />
                    <SPLIT distance="350" swimtime="00:05:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1287" points="326" reactiontime="+84" swimtime="00:03:17.20" resultid="6024" heatid="6181" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:33.55" />
                    <SPLIT distance="150" swimtime="00:02:26.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-25" firstname="Łukasz" gender="M" lastname="Widzik" nation="POL" athleteid="4762">
              <RESULTS>
                <RESULT eventid="1092" points="409" reactiontime="+78" swimtime="00:06:06.21" resultid="4763" heatid="6485" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:21.10" />
                    <SPLIT distance="150" swimtime="00:02:07.04" />
                    <SPLIT distance="200" swimtime="00:02:52.71" />
                    <SPLIT distance="250" swimtime="00:03:44.20" />
                    <SPLIT distance="300" swimtime="00:04:37.70" />
                    <SPLIT distance="350" swimtime="00:05:22.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-02-06" firstname="Dorota" gender="F" lastname="Macoszek" nation="POL" athleteid="4764">
              <RESULTS>
                <RESULT eventid="1595" points="210" reactiontime="+83" swimtime="00:01:58.57" resultid="6501" heatid="6502" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="208" reactiontime="+88" swimtime="00:04:16.17" resultid="4778" heatid="6101" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.13" />
                    <SPLIT distance="100" swimtime="00:01:57.12" />
                    <SPLIT distance="150" swimtime="00:03:05.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="PSK Žilina" nation="SVK">
          <CONTACT name="s" />
          <ATHLETES>
            <ATHLETE birthdate="1960-01-01" firstname="Rastislav" gender="M" lastname="Pavlík" nation="SVK" athleteid="4769">
              <RESULTS>
                <RESULT eventid="1393" status="DNS" swimtime="00:00:00.00" resultid="4770" heatid="6260" lane="6" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Roman" gender="M" lastname="Hrmel" nation="SVK" athleteid="4771">
              <RESULTS>
                <RESULT eventid="1393" points="556" reactiontime="+74" swimtime="00:01:19.10" resultid="4772" heatid="6256" lane="5" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Martin" gender="M" lastname="Strnad" nation="SVK" athleteid="4773">
              <RESULTS>
                <RESULT eventid="1333" points="450" reactiontime="+111" swimtime="00:00:42.00" resultid="4774" heatid="6206" lane="3" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Jaroš" gender="M" lastname="Juraj" nation="SVK" athleteid="4775">
              <RESULTS>
                <RESULT eventid="1333" points="626" swimtime="00:00:37.63" resultid="4776" heatid="6212" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1415" swimtime="00:02:04.25" resultid="4777" heatid="6530" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:06.08" />
                    <SPLIT distance="150" swimtime="00:01:36.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4771" number="1" />
                    <RELAYPOSITION athleteid="4775" number="2" />
                    <RELAYPOSITION athleteid="4769" number="3" />
                    <RELAYPOSITION athleteid="4773" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" name="Azs Uwm Masters Olsztyn" nation="POL">
          <CONTACT city="ŁUPSTYCH" email="gozdzik@uwm.edu.pl" name="Goździejewska Anna" phone="501372846" state="WARM-" street="Leśna1" zip="11-041" />
          <ATHLETES>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="4790">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="4791" heatid="6430" lane="4" />
                <RESULT eventid="1122" points="631" swimtime="00:11:58.86" resultid="4792" heatid="6445" lane="1" entrytime="00:11:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                    <SPLIT distance="100" swimtime="00:01:23.88" />
                    <SPLIT distance="200" swimtime="00:02:58.95" />
                    <SPLIT distance="300" swimtime="00:04:25.05" />
                    <SPLIT distance="400" swimtime="00:05:56.45" />
                    <SPLIT distance="500" swimtime="00:07:27.07" />
                    <SPLIT distance="600" swimtime="00:08:58.15" />
                    <SPLIT distance="700" swimtime="00:10:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="592" reactiontime="+90" swimtime="00:03:23.83" resultid="4793" heatid="6106" lane="5" entrytime="00:03:25.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.51" />
                    <SPLIT distance="100" swimtime="00:01:38.03" />
                    <SPLIT distance="150" swimtime="00:02:30.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="598" reactiontime="+86" swimtime="00:01:15.38" resultid="4794" heatid="6156" lane="5" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="619" reactiontime="+85" swimtime="00:02:41.86" resultid="4795" heatid="6273" lane="5" entrytime="00:03:30.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:19.67" />
                    <SPLIT distance="150" swimtime="00:02:01.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1452" points="592" reactiontime="+80" swimtime="00:03:09.45" resultid="4796" heatid="6296" lane="2" entrytime="00:03:10.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:31.26" />
                    <SPLIT distance="150" swimtime="00:02:24.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="589" reactiontime="+83" swimtime="00:00:33.58" resultid="4797" heatid="6336" lane="2" entrytime="00:00:33.88" />
                <RESULT eventid="1625" points="611" reactiontime="+84" swimtime="00:05:45.19" resultid="4798" heatid="6557" lane="2" entrytime="00:05:42.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:01:22.01" />
                    <SPLIT distance="150" swimtime="00:02:06.22" />
                    <SPLIT distance="200" swimtime="00:02:50.91" />
                    <SPLIT distance="250" swimtime="00:03:35.45" />
                    <SPLIT distance="300" swimtime="00:04:19.77" />
                    <SPLIT distance="350" swimtime="00:05:03.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="4799">
              <RESULTS>
                <RESULT eventid="1092" points="796" reactiontime="+86" swimtime="00:05:41.19" resultid="4800" heatid="6491" lane="3" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:11.96" />
                    <SPLIT distance="150" swimtime="00:01:55.98" />
                    <SPLIT distance="200" swimtime="00:02:39.54" />
                    <SPLIT distance="250" swimtime="00:03:30.86" />
                    <SPLIT distance="300" swimtime="00:04:22.53" />
                    <SPLIT distance="350" swimtime="00:05:03.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="827" reactiontime="+88" swimtime="00:01:09.80" resultid="4801" heatid="6096" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="806" reactiontime="+95" swimtime="00:02:41.39" resultid="4802" heatid="6190" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                    <SPLIT distance="100" swimtime="00:01:18.66" />
                    <SPLIT distance="150" swimtime="00:02:01.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1437" points="787" reactiontime="+92" swimtime="00:02:14.61" resultid="4803" heatid="6289" lane="3" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:06.15" />
                    <SPLIT distance="150" swimtime="00:01:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" points="744" reactiontime="+97" swimtime="00:02:43.89" resultid="4804" heatid="6309" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:07.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="827" reactiontime="+87" swimtime="00:01:07.29" resultid="4805" heatid="6324" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1640" status="DNS" swimtime="00:00:00.00" resultid="4806" heatid="6569" lane="5" entrytime="00:04:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-13" firstname="Michał" gender="M" lastname="Kozikowski" nation="POL" athleteid="4807">
              <RESULTS>
                <RESULT eventid="1228" points="460" reactiontime="+62" swimtime="00:00:33.80" resultid="4808" heatid="6135" lane="2" entrytime="00:00:33.23" />
                <RESULT eventid="1333" points="603" reactiontime="+75" swimtime="00:00:34.87" resultid="4809" heatid="6213" lane="1" entrytime="00:00:36.32" />
                <RESULT comment="O4 - przedwczesny start." eventid="1528" reactiontime="+45" status="DSQ" swimtime="00:00:27.61" resultid="4810" heatid="6351" lane="3" entrytime="00:00:30.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="4811">
              <RESULTS>
                <RESULT eventid="1092" points="540" reactiontime="+84" swimtime="00:05:50.35" resultid="4812" heatid="6491" lane="6" entrytime="00:05:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:16.05" />
                    <SPLIT distance="150" swimtime="00:02:04.56" />
                    <SPLIT distance="200" swimtime="00:02:50.43" />
                    <SPLIT distance="250" swimtime="00:03:41.74" />
                    <SPLIT distance="300" swimtime="00:04:30.03" />
                    <SPLIT distance="350" swimtime="00:05:11.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="596" reactiontime="+83" swimtime="00:01:09.37" resultid="4813" heatid="6096" lane="1" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="632" reactiontime="+53" swimtime="00:00:59.91" resultid="4814" heatid="6172" lane="2" entrytime="00:01:02.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1363" points="675" reactiontime="+81" swimtime="00:00:28.65" resultid="4815" heatid="6237" lane="1" entrytime="00:00:29.93" />
                <RESULT eventid="1467" points="522" reactiontime="+85" swimtime="00:02:35.78" resultid="4816" heatid="6308" lane="6" entrytime="00:02:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:12.72" />
                    <SPLIT distance="150" swimtime="00:01:59.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="663" reactiontime="+79" swimtime="00:00:26.54" resultid="4817" heatid="6360" lane="5" entrytime="00:00:26.90" />
                <RESULT eventid="1610" points="515" reactiontime="+81" swimtime="00:01:18.92" resultid="4818" heatid="6404" lane="1" entrytime="00:01:21.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="AZS Wrocław" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1959-11-21" firstname="Piotr" gender="M" lastname="Figiel" nation="POL" athleteid="6031">
              <RESULTS>
                <RESULT eventid="1168" points="510" reactiontime="+95" swimtime="00:01:21.97" resultid="6032" heatid="6083" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="558" reactiontime="+86" swimtime="00:00:37.19" resultid="6033" heatid="6126" lane="1" />
                <RESULT eventid="1393" points="450" reactiontime="+66" swimtime="00:01:27.65" resultid="6034" heatid="6249" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1467" status="DNS" swimtime="00:00:00.00" resultid="6035" heatid="6299" lane="2" />
                <RESULT eventid="1528" points="494" reactiontime="+100" swimtime="00:00:32.09" resultid="6036" heatid="6341" lane="4" />
                <RESULT eventid="1558" points="359" reactiontime="+78" swimtime="00:03:29.41" resultid="6037" heatid="6372" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:35.17" />
                    <SPLIT distance="150" swimtime="00:02:31.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Michał Derewecki" version="11.75640">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Poznań" name="XXIII Otwarte Integracyjne Mistrzostwa Wielkopolski w Pływaniu w kategoriach Masters" course="SCM" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2023-02-25" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Poznań" nation="POL" />
      <POINTTABLE pointtableid="1126" name="DSV Master Performance Table" version="2022" />
      <QUALIFY from="2021-11-01" until="2023-02-24" />
      <SESSIONS>
        <SESSION date="2023-02-25" daytime="14:55" endtime="19:03" number="1">
          <EVENTS>
            <EVENT eventid="1058" daytime="14:56" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1060" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="1061" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="1062" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7593" />
                    <RANKING order="2" place="2" resultid="7437" />
                    <RANKING order="3" place="3" resultid="7653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7222" />
                    <RANKING order="2" place="2" resultid="7679" />
                    <RANKING order="3" place="3" resultid="7126" />
                    <RANKING order="4" place="4" resultid="7287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7107" />
                    <RANKING order="2" place="2" resultid="7392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7597" />
                    <RANKING order="2" place="2" resultid="7261" />
                    <RANKING order="3" place="3" resultid="7196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7218" />
                    <RANKING order="2" place="2" resultid="7601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="1070" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7562" />
                    <RANKING order="2" place="2" resultid="7151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="1072" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="1073" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="1074" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="1059" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7743" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7744" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" daytime="15:02" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3733" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3734" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3735" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7344" />
                    <RANKING order="2" place="2" resultid="7283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3736" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7690" />
                    <RANKING order="2" place="2" resultid="7364" />
                    <RANKING order="3" place="3" resultid="7116" />
                    <RANKING order="4" place="-1" resultid="7234" />
                    <RANKING order="5" place="-1" resultid="7460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3737" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7181" />
                    <RANKING order="2" place="2" resultid="7675" />
                    <RANKING order="3" place="3" resultid="7238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3738" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7632" />
                    <RANKING order="2" place="2" resultid="7577" />
                    <RANKING order="3" place="3" resultid="7628" />
                    <RANKING order="4" place="4" resultid="7541" />
                    <RANKING order="5" place="5" resultid="7399" />
                    <RANKING order="6" place="6" resultid="7565" />
                    <RANKING order="7" place="7" resultid="7456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3739" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7545" />
                    <RANKING order="2" place="2" resultid="7360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3740" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7573" />
                    <RANKING order="2" place="2" resultid="7205" />
                    <RANKING order="3" place="3" resultid="7395" />
                    <RANKING order="4" place="4" resultid="7252" />
                    <RANKING order="5" place="5" resultid="7581" />
                    <RANKING order="6" place="6" resultid="7604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3741" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7121" />
                    <RANKING order="2" place="2" resultid="7639" />
                    <RANKING order="3" place="-1" resultid="7569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3742" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7452" />
                    <RANKING order="2" place="-1" resultid="7102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3743" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7372" />
                    <RANKING order="2" place="-1" resultid="7585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3744" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3745" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3746" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3747" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3748" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7745" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7746" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7747" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7748" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1093" daytime="15:12" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7026" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="7027" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7028" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="7029" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7536" />
                    <RANKING order="2" place="2" resultid="7654" />
                    <RANKING order="3" place="3" resultid="7438" />
                    <RANKING order="4" place="4" resultid="7130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7030" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7031" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7474" />
                    <RANKING order="2" place="2" resultid="7463" />
                    <RANKING order="3" place="3" resultid="7291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7032" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7598" />
                    <RANKING order="2" place="2" resultid="7471" />
                    <RANKING order="3" place="3" resultid="7403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7033" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7186" />
                    <RANKING order="2" place="2" resultid="7213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7034" agemax="64" agemin="60" name="Kat. H" />
                <AGEGROUP agegroupid="7035" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7036" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7406" />
                    <RANKING order="2" place="2" resultid="7176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7037" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7139" />
                    <RANKING order="2" place="2" resultid="7155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7038" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7265" />
                    <RANKING order="2" place="2" resultid="7162" />
                    <RANKING order="3" place="3" resultid="7159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7039" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="7040" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="7041" agemax="99" agemin="95" name="Kat. O" />
                <AGEGROUP agegroupid="7042" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7608" />
                    <RANKING order="2" place="2" resultid="7536" />
                    <RANKING order="3" place="3" resultid="7186" />
                    <RANKING order="4" place="4" resultid="7598" />
                    <RANKING order="5" place="5" resultid="7654" />
                    <RANKING order="6" place="6" resultid="7471" />
                    <RANKING order="7" place="7" resultid="7438" />
                    <RANKING order="8" place="8" resultid="7474" />
                    <RANKING order="9" place="9" resultid="7463" />
                    <RANKING order="10" place="10" resultid="7213" />
                    <RANKING order="11" place="11" resultid="7403" />
                    <RANKING order="12" place="12" resultid="7130" />
                    <RANKING order="13" place="13" resultid="7406" />
                    <RANKING order="14" place="14" resultid="7291" />
                    <RANKING order="15" place="15" resultid="7549" />
                    <RANKING order="16" place="16" resultid="7265" />
                    <RANKING order="17" place="17" resultid="7467" />
                    <RANKING order="18" place="18" resultid="7176" />
                    <RANKING order="19" place="19" resultid="7139" />
                    <RANKING order="20" place="20" resultid="7162" />
                    <RANKING order="21" place="21" resultid="7155" />
                    <RANKING order="22" place="22" resultid="7159" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7749" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7750" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7751" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1110" daytime="15:20" gender="M" number="4" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3765" agemax="24" agemin="20" name="Kat.0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3766" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3767" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7493" />
                    <RANKING order="2" place="2" resultid="7615" />
                    <RANKING order="3" place="3" resultid="7201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3768" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7117" />
                    <RANKING order="2" place="2" resultid="7349" />
                    <RANKING order="3" place="3" resultid="7279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3769" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7499" />
                    <RANKING order="2" place="2" resultid="7239" />
                    <RANKING order="3" place="3" resultid="7310" />
                    <RANKING order="4" place="-1" resultid="7412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3770" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7588" />
                    <RANKING order="2" place="2" resultid="7301" />
                    <RANKING order="3" place="3" resultid="7425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3771" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7480" />
                    <RANKING order="2" place="2" resultid="7618" />
                    <RANKING order="3" place="3" resultid="7683" />
                    <RANKING order="4" place="4" resultid="7209" />
                    <RANKING order="5" place="5" resultid="7361" />
                    <RANKING order="6" place="6" resultid="7442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3772" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7612" />
                    <RANKING order="2" place="2" resultid="7092" />
                    <RANKING order="3" place="3" resultid="7605" />
                    <RANKING order="4" place="4" resultid="7490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3773" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7409" />
                    <RANKING order="2" place="2" resultid="7387" />
                    <RANKING order="3" place="3" resultid="7483" />
                    <RANKING order="4" place="4" resultid="7486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3774" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3775" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7172" />
                    <RANKING order="2" place="2" resultid="7496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3776" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7477" />
                    <RANKING order="2" place="2" resultid="7447" />
                    <RANKING order="3" place="3" resultid="7143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3777" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3778" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3779" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3780" agemax="99" agemin="95" name="Kat. O" />
                <AGEGROUP agegroupid="6050" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7493" />
                    <RANKING order="2" place="2" resultid="7615" />
                    <RANKING order="3" place="3" resultid="7670" />
                    <RANKING order="4" place="4" resultid="7588" />
                    <RANKING order="5" place="5" resultid="7201" />
                    <RANKING order="6" place="6" resultid="7612" />
                    <RANKING order="7" place="7" resultid="7297" />
                    <RANKING order="8" place="8" resultid="7301" />
                    <RANKING order="9" place="9" resultid="7480" />
                    <RANKING order="10" place="10" resultid="7618" />
                    <RANKING order="11" place="11" resultid="7092" />
                    <RANKING order="12" place="12" resultid="7409" />
                    <RANKING order="13" place="13" resultid="7683" />
                    <RANKING order="14" place="14" resultid="7499" />
                    <RANKING order="15" place="15" resultid="7239" />
                    <RANKING order="16" place="16" resultid="7387" />
                    <RANKING order="17" place="17" resultid="7117" />
                    <RANKING order="18" place="18" resultid="7209" />
                    <RANKING order="19" place="19" resultid="7605" />
                    <RANKING order="20" place="20" resultid="7477" />
                    <RANKING order="21" place="21" resultid="7483" />
                    <RANKING order="22" place="22" resultid="7490" />
                    <RANKING order="23" place="23" resultid="7486" />
                    <RANKING order="24" place="24" resultid="7361" />
                    <RANKING order="25" place="25" resultid="7310" />
                    <RANKING order="26" place="26" resultid="7425" />
                    <RANKING order="27" place="27" resultid="7349" />
                    <RANKING order="28" place="28" resultid="7442" />
                    <RANKING order="29" place="29" resultid="7172" />
                    <RANKING order="30" place="30" resultid="7279" />
                    <RANKING order="31" place="31" resultid="7147" />
                    <RANKING order="32" place="32" resultid="7496" />
                    <RANKING order="33" place="33" resultid="7447" />
                    <RANKING order="34" place="34" resultid="7227" />
                    <RANKING order="35" place="35" resultid="7143" />
                    <RANKING order="36" place="-1" resultid="7412" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7752" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7753" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7754" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7755" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1128" daytime="15:26" gender="F" number="5" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3781" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3782" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="3783" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="3784" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7622" />
                    <RANKING order="2" place="2" resultid="7131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3785" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7193" />
                    <RANKING order="2" place="2" resultid="7506" />
                    <RANKING order="3" place="3" resultid="7288" />
                    <RANKING order="4" place="4" resultid="7468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3786" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7475" />
                    <RANKING order="2" place="2" resultid="7393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3787" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7472" />
                    <RANKING order="2" place="2" resultid="7197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3788" agemax="59" agemin="55" name="Kat. G" />
                <AGEGROUP agegroupid="3789" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3790" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="3791" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="3792" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="3793" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3794" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3795" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3796" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7756" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7757" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1145" daytime="15:30" gender="M" number="6" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3797" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3798" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3799" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7663" />
                    <RANKING order="2" place="2" resultid="7415" />
                    <RANKING order="3" place="3" resultid="7345" />
                    <RANKING order="4" place="4" resultid="7242" />
                    <RANKING order="5" place="5" resultid="7165" />
                    <RANKING order="6" place="6" resultid="7667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3800" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7691" />
                    <RANKING order="2" place="2" resultid="7248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3801" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7182" />
                    <RANKING order="2" place="2" resultid="7676" />
                    <RANKING order="3" place="3" resultid="7082" />
                    <RANKING order="4" place="4" resultid="7078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3802" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7636" />
                    <RANKING order="2" place="2" resultid="7629" />
                    <RANKING order="3" place="3" resultid="7375" />
                    <RANKING order="4" place="4" resultid="7400" />
                    <RANKING order="5" place="5" resultid="7646" />
                    <RANKING order="6" place="6" resultid="7457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3803" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7383" />
                    <RANKING order="2" place="2" resultid="7684" />
                    <RANKING order="3" place="3" resultid="7087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3804" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7574" />
                    <RANKING order="2" place="2" resultid="7253" />
                    <RANKING order="3" place="3" resultid="7582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3805" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7122" />
                    <RANKING order="2" place="-1" resultid="7570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3806" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7230" />
                    <RANKING order="2" place="2" resultid="7111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3807" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="3808" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3809" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3810" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3811" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3812" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7758" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7759" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7760" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1162" daytime="15:36" gender="F" number="7" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3813" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3814" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="3815" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="3816" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7623" />
                    <RANKING order="2" place="-1" resultid="7594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3817" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3818" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7464" />
                    <RANKING order="2" place="2" resultid="7509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3819" agemax="54" agemin="50" name="Kat. F" />
                <AGEGROUP agegroupid="3820" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7512" />
                    <RANKING order="2" place="2" resultid="7602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3821" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3822" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="3823" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7177" />
                    <RANKING order="2" place="2" resultid="7152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3824" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3825" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3826" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3827" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3828" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7761" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7762" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1179" daytime="15:40" gender="M" number="8" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3829" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3830" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="3831" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="3832" agemax="39" agemin="35" name="Kat. C" />
                <AGEGROUP agegroupid="3833" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7427" />
                    <RANKING order="2" place="2" resultid="7336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3834" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7633" />
                    <RANKING order="2" place="2" resultid="7378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3835" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3836" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7396" />
                    <RANKING order="2" place="2" resultid="7093" />
                    <RANKING order="3" place="3" resultid="7271" />
                    <RANKING order="4" place="4" resultid="7367" />
                    <RANKING order="5" place="5" resultid="7275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3837" agemax="64" agemin="60" name="Kat. H" />
                <AGEGROUP agegroupid="3838" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7453" />
                    <RANKING order="2" place="2" resultid="7103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3839" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7527" />
                    <RANKING order="2" place="2" resultid="7552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3840" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7136" />
                    <RANKING order="2" place="2" resultid="7144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3841" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3842" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3843" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3844" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7763" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7764" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1196" daytime="15:46" gender="F" number="9" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3845" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3846" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3847" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3848" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7537" />
                    <RANKING order="2" place="2" resultid="7624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3849" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7127" />
                    <RANKING order="2" place="2" resultid="7507" />
                    <RANKING order="3" place="3" resultid="7680" />
                    <RANKING order="4" place="4" resultid="7469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3850" agemax="49" agemin="45" name="Kat. E" />
                <AGEGROUP agegroupid="3851" agemax="54" agemin="50" name="Kat. F" />
                <AGEGROUP agegroupid="3852" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7187" />
                    <RANKING order="2" place="2" resultid="7513" />
                    <RANKING order="3" place="3" resultid="7214" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3853" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3854" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7169" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3855" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="3856" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7140" />
                    <RANKING order="2" place="2" resultid="7157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3857" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7160" />
                    <RANKING order="2" place="2" resultid="7163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3858" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3859" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3860" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7765" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7766" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1213" daytime="15:50" gender="M" number="10" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3861" agemax="24" agemin="20" name="Kat.0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3862" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="3863" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7664" />
                    <RANKING order="2" place="2" resultid="7346" />
                    <RANKING order="3" place="3" resultid="7243" />
                    <RANKING order="4" place="4" resultid="7202" />
                    <RANKING order="5" place="5" resultid="7166" />
                    <RANKING order="6" place="6" resultid="7245" />
                    <RANKING order="7" place="7" resultid="7668" />
                    <RANKING order="8" place="8" resultid="7284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3864" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7692" />
                    <RANKING order="2" place="2" resultid="7235" />
                    <RANKING order="3" place="3" resultid="7461" />
                    <RANKING order="4" place="4" resultid="7515" />
                    <RANKING order="5" place="5" resultid="7280" />
                    <RANKING order="6" place="6" resultid="7365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3865" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7183" />
                    <RANKING order="2" place="2" resultid="7083" />
                    <RANKING order="3" place="3" resultid="7433" />
                    <RANKING order="4" place="4" resultid="7428" />
                    <RANKING order="5" place="5" resultid="7079" />
                    <RANKING order="6" place="6" resultid="7311" />
                    <RANKING order="7" place="7" resultid="7500" />
                    <RANKING order="8" place="8" resultid="7240" />
                    <RANKING order="9" place="9" resultid="7337" />
                    <RANKING order="10" place="-1" resultid="7413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3866" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7258" />
                    <RANKING order="2" place="2" resultid="7578" />
                    <RANKING order="3" place="3" resultid="7647" />
                    <RANKING order="4" place="4" resultid="7401" />
                    <RANKING order="5" place="5" resultid="7430" />
                    <RANKING order="6" place="6" resultid="7566" />
                    <RANKING order="7" place="7" resultid="7458" />
                    <RANKING order="8" place="8" resultid="7302" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3867" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7546" />
                    <RANKING order="2" place="2" resultid="7210" />
                    <RANKING order="3" place="3" resultid="7619" />
                    <RANKING order="4" place="4" resultid="7362" />
                    <RANKING order="5" place="5" resultid="7088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3868" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7613" />
                    <RANKING order="2" place="2" resultid="7397" />
                    <RANKING order="3" place="3" resultid="7094" />
                    <RANKING order="4" place="4" resultid="7532" />
                    <RANKING order="5" place="5" resultid="7606" />
                    <RANKING order="6" place="6" resultid="7368" />
                    <RANKING order="7" place="7" resultid="7583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3869" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7123" />
                    <RANKING order="2" place="2" resultid="7487" />
                    <RANKING order="3" place="3" resultid="7388" />
                    <RANKING order="4" place="-1" resultid="7571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3870" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7231" />
                    <RANKING order="2" place="2" resultid="7686" />
                    <RANKING order="3" place="3" resultid="7112" />
                    <RANKING order="4" place="4" resultid="7148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3871" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7528" />
                    <RANKING order="2" place="2" resultid="7173" />
                    <RANKING order="3" place="3" resultid="7373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3872" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7098" />
                    <RANKING order="2" place="2" resultid="7448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3873" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3874" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3875" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3876" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7767" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7768" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7769" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7770" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7771" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7772" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7044" daytime="15:58" gender="F" number="11" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7045" agemax="99" agemin="80" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="7046" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL" />
                <AGEGROUP agegroupid="7047" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL" />
                <AGEGROUP agegroupid="7048" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL" />
                <AGEGROUP agegroupid="7049" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7050" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL" />
                <AGEGROUP agegroupid="7051" agemax="400" agemin="280" name="Kat. F" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7773" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1247" daytime="16:04" gender="M" number="12" order="13" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4005" agemax="99" agemin="80" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="4006" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL" />
                <AGEGROUP agegroupid="4007" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4008" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7522" />
                    <RANKING order="2" place="2" resultid="7434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4009" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7625" />
                    <RANKING order="2" place="2" resultid="7523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4010" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL" />
                <AGEGROUP agegroupid="4011" agemax="400" agemin="280" name="Kat. F" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7774" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7052" daytime="16:10" gender="X" number="13" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7053" agemax="99" agemin="80" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="7054" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL" />
                <AGEGROUP agegroupid="7055" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL" />
                <AGEGROUP agegroupid="7056" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7626" />
                    <RANKING order="2" place="-1" resultid="7422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7057" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7524" />
                    <RANKING order="2" place="2" resultid="7293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7058" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7059" agemax="400" agemin="280" name="Kat. F" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7775" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7068" daytime="16:20" gender="F" number="14" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7069" agemax="-1" agemin="1" name="Niepełnosprawni">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7314" />
                    <RANKING order="2" place="2" resultid="7318" />
                    <RANKING order="3" place="3" resultid="7316" />
                    <RANKING order="4" place="4" resultid="7320" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7776" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1298" daytime="16:22" gender="M" number="15" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1332" agemax="-1" agemin="1" name="Niepełnosprawni">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7685" />
                    <RANKING order="2" place="2" resultid="7341" />
                    <RANKING order="3" place="3" resultid="7322" />
                    <RANKING order="4" place="4" resultid="7326" />
                    <RANKING order="5" place="5" resultid="7328" />
                    <RANKING order="6" place="6" resultid="7324" />
                    <RANKING order="7" place="7" resultid="7338" />
                    <RANKING order="8" place="8" resultid="7269" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7777" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1315" daytime="16:26" gender="F" number="16" order="21" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3877" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3878" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3879" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="3880" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7538" />
                    <RANKING order="2" place="2" resultid="7439" />
                    <RANKING order="3" place="3" resultid="7132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3881" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3882" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7465" />
                    <RANKING order="2" place="2" resultid="7518" />
                    <RANKING order="3" place="3" resultid="7292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3883" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7599" />
                    <RANKING order="2" place="2" resultid="7404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3884" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3885" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3886" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3887" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7407" />
                    <RANKING order="2" place="2" resultid="7178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3888" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="3889" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3890" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3891" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3892" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7778" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7779" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1333" daytime="16:38" gender="M" number="17" order="22" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3893" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3894" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="3895" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7494" />
                    <RANKING order="2" place="2" resultid="7203" />
                    <RANKING order="3" place="3" resultid="7167" />
                    <RANKING order="4" place="4" resultid="7285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3896" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7118" />
                    <RANKING order="2" place="2" resultid="7350" />
                    <RANKING order="3" place="3" resultid="7281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3897" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3898" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7589" />
                    <RANKING order="2" place="2" resultid="7303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3899" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3900" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3901" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7410" />
                    <RANKING order="2" place="2" resultid="7389" />
                    <RANKING order="3" place="3" resultid="7488" />
                    <RANKING order="4" place="4" resultid="7484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3902" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7454" />
                    <RANKING order="2" place="2" resultid="7149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3903" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3904" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7478" />
                    <RANKING order="2" place="2" resultid="7145" />
                    <RANKING order="3" place="-1" resultid="7449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3905" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3906" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3907" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3908" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7780" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7781" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7782" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1350" daytime="16:54" gender="F" number="18" order="23" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3909" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3910" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="3911" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="3912" agemax="39" agemin="35" name="Kat. C" />
                <AGEGROUP agegroupid="3913" agemax="44" agemin="40" name="Kat. D" />
                <AGEGROUP agegroupid="3914" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3915" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3916" agemax="59" agemin="55" name="Kat. G" />
                <AGEGROUP agegroupid="3917" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7191" />
                    <RANKING order="2" place="2" resultid="7557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3918" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="3919" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="3920" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="3921" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3922" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3923" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3924" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7783" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1367" daytime="17:00" gender="M" number="19" order="24" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3925" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3926" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3927" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="3928" agemax="39" agemin="35" name="Kat. C" />
                <AGEGROUP agegroupid="3929" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7420" />
                    <RANKING order="2" place="-1" resultid="7677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3930" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7542" />
                    <RANKING order="2" place="2" resultid="7630" />
                    <RANKING order="3" place="3" resultid="7376" />
                    <RANKING order="4" place="-1" resultid="7648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3931" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3932" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7272" />
                    <RANKING order="2" place="2" resultid="7491" />
                    <RANKING order="3" place="3" resultid="7276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3933" agemax="64" agemin="60" name="Kat. H" />
                <AGEGROUP agegroupid="3934" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="3935" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="3936" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="3937" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3938" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3939" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3940" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7784" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7785" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1384" daytime="17:10" gender="F" number="20" order="25" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3941" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3942" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="3943" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3944" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3945" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7223" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3946" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3947" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7262" />
                    <RANKING order="2" place="2" resultid="7198" />
                    <RANKING order="3" place="3" resultid="7332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3948" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7188" />
                    <RANKING order="2" place="2" resultid="7219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3949" agemax="64" agemin="60" name="Kat. H" />
                <AGEGROUP agegroupid="3950" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3951" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3952" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3953" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3954" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3955" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3956" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7786" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7787" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1401" daytime="17:24" gender="M" number="21" order="26" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3957" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3958" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="3959" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="3960" agemax="39" agemin="35" name="Kat. C" />
                <AGEGROUP agegroupid="3961" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3962" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7637" />
                    <RANKING order="2" place="2" resultid="7634" />
                    <RANKING order="3" place="3" resultid="7379" />
                    <RANKING order="4" place="-1" resultid="7431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3963" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7384" />
                    <RANKING order="2" place="2" resultid="7547" />
                    <RANKING order="3" place="3" resultid="7444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3964" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7575" />
                    <RANKING order="2" place="2" resultid="7273" />
                    <RANKING order="3" place="3" resultid="7369" />
                    <RANKING order="4" place="4" resultid="7277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3965" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3966" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3967" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7586" />
                    <RANKING order="2" place="-1" resultid="7553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3968" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3969" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3970" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3971" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3972" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7788" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7789" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1418" daytime="17:34" gender="F" number="22" order="27" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3973" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3974" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="3975" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="3976" agemax="39" agemin="35" name="Kat. C" />
                <AGEGROUP agegroupid="3977" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7224" />
                    <RANKING order="2" place="2" resultid="7128" />
                    <RANKING order="3" place="3" resultid="7681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3978" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7108" />
                    <RANKING order="2" place="2" resultid="7520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3979" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3980" agemax="59" agemin="55" name="Kat. G" />
                <AGEGROUP agegroupid="3981" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7558" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3982" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="3983" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3984" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="3985" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="3986" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="3987" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="3988" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7790" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1435" daytime="17:54" gender="M" number="23" order="28" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3989" agemax="24" agemin="20" name="Kat.0" />
                <AGEGROUP agegroupid="3990" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="3991" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7616" />
                    <RANKING order="2" place="2" resultid="7246" />
                    <RANKING order="3" place="3" resultid="7416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3992" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7249" />
                    <RANKING order="2" place="-1" resultid="7793" />
                    <RANKING order="3" place="-1" resultid="7516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3993" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3994" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7579" />
                    <RANKING order="2" place="2" resultid="7590" />
                    <RANKING order="3" place="3" resultid="7567" />
                    <RANKING order="4" place="4" resultid="7380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3995" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3996" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7206" />
                    <RANKING order="2" place="2" resultid="7651" />
                    <RANKING order="3" place="-1" resultid="7533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3997" agemax="64" agemin="60" name="Kat. H" />
                <AGEGROUP agegroupid="3998" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3999" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7529" />
                    <RANKING order="2" place="2" resultid="7554" />
                    <RANKING order="3" place="3" resultid="7174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4000" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4001" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="4002" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="4003" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="4004" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7791" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7792" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="7390" name="KS Warta Poznań">
          <ATHLETES>
            <ATHLETE firstname="Błażej" lastname="Wachowski" birthdate="1980-10-08" gender="M" nation="POL" license="100115700545" swrid="4595659" athleteid="7419">
              <RESULTS>
                <RESULT eventid="1367" points="465" reactiontime="+77" swimtime="00:02:42.65" resultid="7420" heatid="7785" lane="6" entrytime="00:02:38.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="150" swimtime="00:02:00.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="514" swimtime="00:10:38.53" resultid="7421" heatid="7792" lane="2" entrytime="00:10:20.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:14.88" />
                    <SPLIT distance="150" swimtime="00:01:54.86" />
                    <SPLIT distance="200" swimtime="00:02:35.09" />
                    <SPLIT distance="250" swimtime="00:03:15.45" />
                    <SPLIT distance="300" swimtime="00:03:55.92" />
                    <SPLIT distance="350" swimtime="00:04:36.61" />
                    <SPLIT distance="400" swimtime="00:05:17.44" />
                    <SPLIT distance="450" swimtime="00:05:57.73" />
                    <SPLIT distance="500" swimtime="00:06:38.43" />
                    <SPLIT distance="550" swimtime="00:07:19.24" />
                    <SPLIT distance="600" swimtime="00:08:00.20" />
                    <SPLIT distance="650" swimtime="00:08:40.82" />
                    <SPLIT distance="700" swimtime="00:09:21.52" />
                    <SPLIT distance="750" swimtime="00:10:01.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Janyga" birthdate="1966-03-27" gender="M" nation="POL" license="100115700346" swrid="4992782" athleteid="7394">
              <RESULTS>
                <RESULT eventid="1075" points="782" reactiontime="+71" swimtime="00:01:11.34" resultid="7395" heatid="7748" lane="0" entrytime="00:01:11.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="674" reactiontime="+69" swimtime="00:00:33.46" resultid="7396" heatid="7764" lane="5" entrytime="00:00:32.07" entrycourse="SCM" />
                <RESULT eventid="1213" points="737" reactiontime="+71" swimtime="00:00:28.81" resultid="7397" heatid="7771" lane="3" entrytime="00:00:28.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Zawadka" birthdate="1978-12-30" gender="M" nation="POL" license="500115700748" athleteid="7398">
              <RESULTS>
                <RESULT eventid="1075" points="507" reactiontime="+85" swimtime="00:01:15.22" resultid="7399" heatid="7747" lane="3" entrytime="00:01:16.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="527" reactiontime="+80" swimtime="00:00:31.78" resultid="7400" heatid="7758" lane="3" entrytime="00:00:33.26" />
                <RESULT eventid="1213" points="492" reactiontime="+74" swimtime="00:00:30.22" resultid="7401" heatid="7770" lane="1" entrytime="00:00:31.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Kuca" birthdate="1994-07-23" gender="M" nation="POL" license="100115700396" swrid="4213120" athleteid="7417">
              <RESULTS>
                <RESULT eventid="1367" points="954" swimtime="00:02:08.25" resultid="7418" heatid="7785" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                    <SPLIT distance="100" swimtime="00:00:59.55" />
                    <SPLIT distance="150" swimtime="00:01:33.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Waraczewski" birthdate="1962-04-19" gender="M" nation="POL" license="100115700344" swrid="4992781" athleteid="7408">
              <RESULTS>
                <RESULT eventid="1110" points="572" swimtime="00:00:39.42" resultid="7409" heatid="7754" lane="4" entrytime="00:00:38.55" entrycourse="SCM" />
                <RESULT eventid="1333" points="688" reactiontime="+98" swimtime="00:03:07.87" resultid="7410" heatid="7782" lane="7" entrytime="00:03:09.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                    <SPLIT distance="100" swimtime="00:01:29.44" />
                    <SPLIT distance="150" swimtime="00:02:18.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szymkowiak" birthdate="1980-04-12" gender="M" nation="POL" license="500115700523" swrid="5312534" athleteid="7411">
              <RESULTS>
                <RESULT eventid="1110" status="DNS" swimtime="00:00:00.00" resultid="7412" heatid="7755" lane="3" entrytime="00:00:30.39" entrycourse="SCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="7413" heatid="7772" lane="6" entrytime="00:00:25.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Krupińska" birthdate="1953-05-24" gender="F" nation="POL" license="500115600520" swrid="4992790" athleteid="7405">
              <RESULTS>
                <RESULT eventid="1093" points="524" swimtime="00:00:53.55" resultid="7406" heatid="7750" lane="4" entrytime="00:00:53.25" entrycourse="SCM" />
                <RESULT eventid="1315" points="592" swimtime="00:04:13.80" resultid="7407" heatid="7778" lane="4" entrytime="00:04:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.42" />
                    <SPLIT distance="100" swimtime="00:02:04.48" />
                    <SPLIT distance="150" swimtime="00:03:11.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sylwia" lastname="Gorockiewicz" birthdate="1975-03-29" gender="F" nation="POL" license="500115600525" swrid="4837788" athleteid="7391">
              <RESULTS>
                <RESULT eventid="1058" points="136" reactiontime="+116" swimtime="00:02:14.28" resultid="7392" heatid="7743" lane="6" entrytime="00:02:13.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="95" reactiontime="+111" swimtime="00:01:05.76" resultid="7393" heatid="7756" lane="5" entrytime="00:01:09.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Witt" birthdate="1991-08-11" gender="M" nation="POL" license="500115700645" swrid="5062813" athleteid="7414">
              <RESULTS>
                <RESULT eventid="1145" points="604" reactiontime="+68" swimtime="00:00:27.05" resultid="7415" heatid="7760" lane="3" entrytime="00:00:26.35" entrycourse="SCM" />
                <RESULT eventid="1435" points="584" reactiontime="+76" swimtime="00:09:56.99" resultid="7416" heatid="7792" lane="3" entrytime="00:09:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="100" swimtime="00:01:06.55" />
                    <SPLIT distance="150" swimtime="00:01:42.88" />
                    <SPLIT distance="200" swimtime="00:02:19.08" />
                    <SPLIT distance="250" swimtime="00:02:55.73" />
                    <SPLIT distance="300" swimtime="00:03:32.73" />
                    <SPLIT distance="350" swimtime="00:04:10.00" />
                    <SPLIT distance="400" swimtime="00:04:47.93" />
                    <SPLIT distance="450" swimtime="00:05:26.40" />
                    <SPLIT distance="500" swimtime="00:06:05.46" />
                    <SPLIT distance="550" swimtime="00:06:43.77" />
                    <SPLIT distance="600" swimtime="00:07:22.83" />
                    <SPLIT distance="650" swimtime="00:08:02.27" />
                    <SPLIT distance="700" swimtime="00:08:41.93" />
                    <SPLIT distance="750" swimtime="00:09:20.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Skurczyńska" birthdate="1971-10-13" gender="F" nation="POL" license="500115600746" athleteid="7402">
              <RESULTS>
                <RESULT eventid="1093" points="401" swimtime="00:00:48.55" resultid="7403" heatid="7751" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="1315" points="355" swimtime="00:03:57.56" resultid="7404" heatid="7779" lane="9" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.91" />
                    <SPLIT distance="100" swimtime="00:01:52.52" />
                    <SPLIT distance="150" swimtime="00:02:57.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="7052" status="DNS" swimtime="00:00:00.00" resultid="7422" heatid="7775" lane="5" entrytime="00:06:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7398" number="1" />
                    <RELAYPOSITION athleteid="7402" number="2" />
                    <RELAYPOSITION athleteid="7411" number="3" />
                    <RELAYPOSITION athleteid="7391" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7217" name="MKP Szczecin">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Serbin" birthdate="1966-01-01" gender="F" nation="POL" swrid="4302596" athleteid="7216">
              <RESULTS>
                <RESULT eventid="1058" points="606" reactiontime="+76" swimtime="00:01:26.18" resultid="7218" heatid="7744" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="656" reactiontime="+75" swimtime="00:03:00.67" resultid="7219" heatid="7787" lane="5" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:01:28.37" />
                    <SPLIT distance="150" swimtime="00:02:15.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7200" name="Start Poznań">
          <ATHLETES>
            <ATHLETE firstname="Zbigniew" lastname="Wróbel" birthdate="1967-01-01" gender="M" nation="POL" athleteid="7251">
              <RESULTS>
                <RESULT eventid="1075" points="777" reactiontime="+90" swimtime="00:01:11.50" resultid="7252" heatid="7748" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="763" reactiontime="+85" swimtime="00:00:30.69" resultid="7253" heatid="7759" lane="5" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Jędrychowski" birthdate="1989-01-01" gender="M" nation="POL" swrid="4285568" athleteid="7199">
              <RESULTS>
                <RESULT eventid="1110" points="644" reactiontime="+73" swimtime="00:00:32.19" resultid="7201" heatid="7755" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1213" points="540" swimtime="00:00:27.17" resultid="7202" heatid="7772" lane="8" entrytime="00:00:27.00" />
                <RESULT eventid="1333" points="638" reactiontime="+83" swimtime="00:02:43.20" resultid="7203" heatid="7782" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:19.27" />
                    <SPLIT distance="150" swimtime="00:02:02.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Monczak" birthdate="1967-01-01" gender="M" nation="POL" swrid="4302571" athleteid="7204">
              <RESULTS>
                <RESULT eventid="1075" points="826" swimtime="00:01:10.06" resultid="7205" heatid="7748" lane="2" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="741" reactiontime="+76" swimtime="00:10:16.58" resultid="7206" heatid="7792" lane="6" entrytime="00:10:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:11.94" />
                    <SPLIT distance="150" swimtime="00:01:50.05" />
                    <SPLIT distance="200" swimtime="00:02:28.36" />
                    <SPLIT distance="250" swimtime="00:03:06.94" />
                    <SPLIT distance="300" swimtime="00:03:45.57" />
                    <SPLIT distance="350" swimtime="00:04:24.40" />
                    <SPLIT distance="400" swimtime="00:05:03.19" />
                    <SPLIT distance="450" swimtime="00:05:41.81" />
                    <SPLIT distance="500" swimtime="00:06:21.32" />
                    <SPLIT distance="550" swimtime="00:07:00.74" />
                    <SPLIT distance="600" swimtime="00:07:40.37" />
                    <SPLIT distance="650" swimtime="00:08:19.75" />
                    <SPLIT distance="700" swimtime="00:08:59.10" />
                    <SPLIT distance="750" swimtime="00:09:38.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7689" name="Masters Lublin">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Dawidek" birthdate="1986-01-01" gender="M" nation="POL" athleteid="7688">
              <RESULTS>
                <RESULT eventid="1075" points="510" reactiontime="+77" swimtime="00:01:11.06" resultid="7690" heatid="7747" lane="5" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="470" reactiontime="+73" swimtime="00:00:30.38" resultid="7691" heatid="7759" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1213" points="509" reactiontime="+74" swimtime="00:00:27.59" resultid="7692" heatid="7772" lane="0" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7295" name="niezrzeszony Poznań">
          <ATHLETES>
            <ATHLETE firstname="Filip" lastname="Wiatrowski" birthdate="1996-01-01" gender="M" nation="POL" swrid="4290292" athleteid="7294">
              <RESULTS>
                <RESULT eventid="1075" points="514" reactiontime="+75" swimtime="00:01:08.91" resultid="7296" heatid="7748" lane="3" entrytime="00:01:07.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1110" points="504" reactiontime="+76" swimtime="00:00:35.51" resultid="7297" heatid="7755" lane="8" entrytime="00:00:34.09" />
                <RESULT eventid="1145" points="452" swimtime="00:00:30.88" resultid="7298" heatid="7760" lane="9" entrytime="00:00:29.13" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="15" clubid="7423" name="KU AZS UAM Poznań">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Juszkiewicz" birthdate="1974-05-10" gender="M" nation="POL" license="503315700077" swrid="5537971" athleteid="7429">
              <RESULTS>
                <RESULT eventid="1213" points="467" reactiontime="+78" swimtime="00:00:30.76" resultid="7430" heatid="7770" lane="3" entrytime="00:00:30.97" entrycourse="SCM" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="7431" heatid="7788" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Strzelczyk" birthdate="1978-07-20" gender="M" nation="POL" license="503315700084" athleteid="7424">
              <RESULTS>
                <RESULT eventid="1110" points="297" swimtime="00:00:45.38" resultid="7425" heatid="7752" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Kaczmarek" birthdate="1983-07-27" gender="M" nation="POL" license="503315700216" swrid="5537972" athleteid="7426">
              <RESULTS>
                <RESULT eventid="1179" points="534" reactiontime="+71" swimtime="00:00:33.46" resultid="7427" heatid="7764" lane="3" entrytime="00:00:33.11" entrycourse="SCM" />
                <RESULT eventid="1213" points="551" reactiontime="+68" swimtime="00:00:28.31" resultid="7428" heatid="7771" lane="6" entrytime="00:00:28.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kaczmarek" birthdate="1982-10-03" gender="M" nation="POL" license="503315700221" swrid="5471723" athleteid="7432">
              <RESULTS>
                <RESULT eventid="1213" points="564" reactiontime="+95" swimtime="00:00:28.08" resultid="7433" heatid="7767" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1247" reactiontime="+71" swimtime="00:05:31.52" resultid="7434" heatid="7774" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:17.26" />
                    <SPLIT distance="150" swimtime="00:02:04.75" />
                    <SPLIT distance="200" swimtime="00:03:01.63" />
                    <SPLIT distance="250" swimtime="00:03:38.13" />
                    <SPLIT distance="300" swimtime="00:04:20.21" />
                    <SPLIT distance="350" swimtime="00:04:54.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7426" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="7424" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="7432" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="7429" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02202" nation="POL" region="02" clubid="7440" name="MKS ,,Astoria&apos;&apos; Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-13" gender="M" nation="POL" license="102202700126" swrid="5471726" athleteid="7441">
              <RESULTS>
                <RESULT eventid="1110" points="273" swimtime="00:00:47.39" resultid="7442" heatid="7753" lane="8" entrytime="00:00:48.74" entrycourse="SCM" />
                <RESULT eventid="1179" points="128" reactiontime="+90" swimtime="00:00:56.15" resultid="7443" heatid="7763" lane="3" entrytime="00:00:53.09" entrycourse="SCM" />
                <RESULT eventid="1401" points="140" reactiontime="+96" swimtime="00:04:27.68" resultid="7444" heatid="7788" lane="3" entrytime="00:04:21.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.40" />
                    <SPLIT distance="150" swimtime="00:03:17.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LARISW" nation="POL" clubid="7347" name="Lubuska Akademia Ratownictwa I Sportów Wodnych">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Krupiński" birthdate="1987-02-05" gender="M" nation="POL" license="501404700235" swrid="5568771" athleteid="7348">
              <RESULTS>
                <RESULT eventid="1110" points="238" reactiontime="+95" swimtime="00:00:46.55" resultid="7349" heatid="7753" lane="7" entrytime="00:00:45.85" />
                <RESULT eventid="1333" points="268" reactiontime="+99" swimtime="00:03:37.89" resultid="7350" heatid="7781" lane="5" entrytime="00:03:35.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.81" />
                    <SPLIT distance="100" swimtime="00:01:44.10" />
                    <SPLIT distance="150" swimtime="00:02:41.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7086" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Łopuszyński" birthdate="1969-01-01" gender="M" nation="POL" athleteid="7085">
              <RESULTS>
                <RESULT eventid="1145" points="177" reactiontime="+108" swimtime="00:00:47.68" resultid="7087" heatid="7758" lane="1" entrytime="00:00:48.00" />
                <RESULT eventid="1213" points="189" swimtime="00:00:42.64" resultid="7088" heatid="7768" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="1367" points="211" reactiontime="+108" swimtime="00:03:53.28" resultid="7089" heatid="7784" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.29" />
                    <SPLIT distance="100" swimtime="00:01:50.29" />
                    <SPLIT distance="150" swimtime="00:02:51.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7091" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Lewandowski" birthdate="1968-01-01" gender="M" nation="POL" swrid="4992668" athleteid="7090">
              <RESULTS>
                <RESULT eventid="1110" points="471" swimtime="00:00:39.19" resultid="7092" heatid="7755" lane="9" entrytime="00:00:38.50" />
                <RESULT eventid="1179" points="336" reactiontime="+77" swimtime="00:00:42.20" resultid="7093" heatid="7764" lane="7" entrytime="00:00:42.20" />
                <RESULT eventid="1213" points="461" swimtime="00:00:33.69" resultid="7094" heatid="7769" lane="4" entrytime="00:00:32.20" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="GBR" clubid="7081" name="Wantage White Horses">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Rybak" birthdate="1980-01-01" gender="M" nation="GBR" athleteid="7080">
              <RESULTS>
                <RESULT eventid="1145" points="656" reactiontime="+80" swimtime="00:00:28.92" resultid="7082" heatid="7760" lane="7" entrytime="00:00:28.62" />
                <RESULT eventid="1213" points="619" reactiontime="+78" swimtime="00:00:27.23" resultid="7083" heatid="7772" lane="7" entrytime="00:00:26.76" />
                <RESULT eventid="1401" points="518" reactiontime="+68" swimtime="00:02:42.41" resultid="7084" heatid="7789" lane="3" entrytime="00:02:50.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:17.25" />
                    <SPLIT distance="150" swimtime="00:01:59.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01203" nation="POL" region="03" clubid="7539" name="UKS ,,Trójka&apos;&apos; Puławy">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Gogacz" birthdate="1976-10-28" gender="M" nation="POL" license="501203700057" swrid="4754646" athleteid="7540">
              <RESULTS>
                <RESULT eventid="1075" points="549" reactiontime="+79" swimtime="00:01:13.25" resultid="7541" heatid="7746" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="607" reactiontime="+79" swimtime="00:02:35.49" resultid="7542" heatid="7785" lane="5" entrytime="00:02:29.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:14.84" />
                    <SPLIT distance="150" swimtime="00:01:55.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7304" name="T.P. Masters Opole" />
        <CLUB type="CLUB" code="03415" nation="POL" region="15" clubid="7543" name="Uks Cityzen">
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Matyszczak" birthdate="1970-12-14" gender="M" nation="POL" license="503415700353" swrid="5471729" athleteid="7544">
              <RESULTS>
                <RESULT eventid="1075" points="357" reactiontime="+90" swimtime="00:01:23.60" resultid="7545" heatid="7747" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="503" reactiontime="+83" swimtime="00:00:30.78" resultid="7546" heatid="7770" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1401" points="322" reactiontime="+85" swimtime="00:03:22.98" resultid="7547" heatid="7789" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rusłana" lastname="Dembecka" birthdate="1957-10-01" gender="F" nation="POL" license="503415600404" athleteid="7548">
              <RESULTS>
                <RESULT eventid="1093" points="333" swimtime="00:00:56.08" resultid="7549" heatid="7750" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="1315" points="403" reactiontime="+119" swimtime="00:04:31.85" resultid="7550" heatid="7778" lane="3" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.11" />
                    <SPLIT distance="100" swimtime="00:02:13.31" />
                    <SPLIT distance="150" swimtime="00:03:23.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Putowska" birthdate="1962-01-22" gender="F" nation="POL" license="503415600402" swrid="5416834" athleteid="7555">
              <RESULTS>
                <RESULT eventid="1315" points="452" swimtime="00:04:04.08" resultid="7556" heatid="7779" lane="0" entrytime="00:03:57.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.20" />
                    <SPLIT distance="100" swimtime="00:01:56.50" />
                    <SPLIT distance="150" swimtime="00:03:00.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="378" swimtime="00:04:40.90" resultid="7557" heatid="7783" lane="6" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.50" />
                    <SPLIT distance="100" swimtime="00:02:11.60" />
                    <SPLIT distance="150" swimtime="00:03:27.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="380" swimtime="00:15:54.94" resultid="7558" heatid="7790" lane="1" entrytime="00:15:39.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.99" />
                    <SPLIT distance="100" swimtime="00:01:47.31" />
                    <SPLIT distance="150" swimtime="00:02:46.76" />
                    <SPLIT distance="200" swimtime="00:03:46.35" />
                    <SPLIT distance="250" swimtime="00:04:46.62" />
                    <SPLIT distance="300" swimtime="00:05:47.72" />
                    <SPLIT distance="350" swimtime="00:06:49.02" />
                    <SPLIT distance="400" swimtime="00:07:49.63" />
                    <SPLIT distance="450" swimtime="00:08:51.37" />
                    <SPLIT distance="500" swimtime="00:09:52.45" />
                    <SPLIT distance="550" swimtime="00:10:53.73" />
                    <SPLIT distance="600" swimtime="00:11:54.10" />
                    <SPLIT distance="650" swimtime="00:12:54.78" />
                    <SPLIT distance="700" swimtime="00:13:56.19" />
                    <SPLIT distance="750" swimtime="00:14:57.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Boryski" birthdate="1951-03-05" gender="M" nation="POL" license="503415700180" swrid="4754708" athleteid="7551">
              <RESULTS>
                <RESULT eventid="1179" points="387" reactiontime="+89" swimtime="00:00:47.58" resultid="7552" heatid="7763" lane="4" entrytime="00:00:48.04" entrycourse="SCM" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="7553" heatid="7788" lane="4" entrytime="00:03:50.88" entrycourse="SCM" />
                <RESULT eventid="1435" points="469" reactiontime="+108" swimtime="00:14:45.43" resultid="7554" heatid="7791" lane="7" entrytime="00:14:53.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                    <SPLIT distance="100" swimtime="00:01:45.19" />
                    <SPLIT distance="150" swimtime="00:02:41.57" />
                    <SPLIT distance="200" swimtime="00:03:37.31" />
                    <SPLIT distance="250" swimtime="00:04:32.83" />
                    <SPLIT distance="300" swimtime="00:05:28.57" />
                    <SPLIT distance="350" swimtime="00:06:24.38" />
                    <SPLIT distance="400" swimtime="00:07:20.57" />
                    <SPLIT distance="450" swimtime="00:08:15.72" />
                    <SPLIT distance="500" swimtime="00:09:11.54" />
                    <SPLIT distance="550" swimtime="00:10:07.51" />
                    <SPLIT distance="600" swimtime="00:11:03.87" />
                    <SPLIT distance="650" swimtime="00:11:59.60" />
                    <SPLIT distance="700" swimtime="00:12:55.25" />
                    <SPLIT distance="750" swimtime="00:13:51.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="7052" reactiontime="+45" swimtime="00:07:10.81" resultid="7559" heatid="7775" lane="3" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.55" />
                    <SPLIT distance="100" swimtime="00:01:48.39" />
                    <SPLIT distance="150" swimtime="00:02:51.22" />
                    <SPLIT distance="200" swimtime="00:03:58.19" />
                    <SPLIT distance="250" swimtime="00:04:52.80" />
                    <SPLIT distance="300" swimtime="00:05:58.75" />
                    <SPLIT distance="350" swimtime="00:06:32.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7551" number="1" reactiontime="+45" />
                    <RELAYPOSITION athleteid="7548" number="2" reactiontime="+104" />
                    <RELAYPOSITION athleteid="7555" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="7544" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7672" name="Niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Wilk" birthdate="1991-01-01" gender="M" nation="POL" athleteid="7665">
              <RESULTS>
                <RESULT eventid="1145" points="415" swimtime="00:00:30.66" resultid="7667" heatid="7759" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1213" points="458" swimtime="00:00:28.69" resultid="7668" heatid="7771" lane="9" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="14814" nation="POL" region="14" clubid="7525" name="Stowarzyszenie Pływackie Legia Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Bogdan" lastname="Dubiński" birthdate="1953-05-05" gender="M" nation="POL" license="514814700003" swrid="4992696" athleteid="7526">
              <RESULTS>
                <RESULT eventid="1179" points="462" reactiontime="+86" swimtime="00:00:44.83" resultid="7527" heatid="7764" lane="1" entrytime="00:00:42.82" entrycourse="SCM" />
                <RESULT eventid="1213" points="532" swimtime="00:00:35.04" resultid="7528" heatid="7768" lane="4" entrytime="00:00:36.23" entrycourse="SCM" />
                <RESULT eventid="1435" points="517" swimtime="00:14:17.02" resultid="7529" heatid="7791" lane="1" entrytime="00:15:34.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:01:34.23" />
                    <SPLIT distance="150" swimtime="00:02:28.16" />
                    <SPLIT distance="200" swimtime="00:03:23.34" />
                    <SPLIT distance="250" swimtime="00:04:17.19" />
                    <SPLIT distance="300" swimtime="00:05:12.81" />
                    <SPLIT distance="350" swimtime="00:06:08.64" />
                    <SPLIT distance="400" swimtime="00:07:04.25" />
                    <SPLIT distance="450" swimtime="00:07:59.67" />
                    <SPLIT distance="500" swimtime="00:08:55.03" />
                    <SPLIT distance="550" swimtime="00:09:50.96" />
                    <SPLIT distance="600" swimtime="00:10:46.13" />
                    <SPLIT distance="650" swimtime="00:11:41.22" />
                    <SPLIT distance="700" swimtime="00:12:35.81" />
                    <SPLIT distance="750" swimtime="00:13:29.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7100" name="UKS SP8 Chrzanów">
          <ATHLETES>
            <ATHLETE firstname="Alfred" lastname="Zabrzański" birthdate="1954-05-12" gender="M" nation="POL" swrid="4477631" athleteid="7101">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="7102" heatid="7747" lane="9" entrytime="00:01:32.00" />
                <RESULT eventid="1179" points="442" reactiontime="+90" swimtime="00:00:43.73" resultid="7103" heatid="7764" lane="8" entrytime="00:00:44.70" />
                <RESULT eventid="1213" points="567" swimtime="00:00:33.32" resultid="7686" heatid="7769" lane="9" entrytime="00:00:34.78" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00607" nation="POL" region="07" clubid="7530" name="Towarzystwo Pływackie ,,Masters&apos;&apos; Opole">
          <ATHLETES>
            <ATHLETE firstname="Grzegorz" lastname="Mandziuk" birthdate="1965-04-11" gender="M" nation="POL" license="100607700033" athleteid="7531">
              <RESULTS>
                <RESULT eventid="1213" points="391" reactiontime="+76" swimtime="00:00:35.57" resultid="7532" heatid="7769" lane="0" entrytime="00:00:34.70" />
                <RESULT eventid="1435" status="OTL" swimtime="00:16:04.80" resultid="7533" heatid="7791" lane="6" entrytime="00:14:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                    <SPLIT distance="100" swimtime="00:01:41.88" />
                    <SPLIT distance="150" swimtime="00:02:42.97" />
                    <SPLIT distance="200" swimtime="00:03:44.47" />
                    <SPLIT distance="250" swimtime="00:04:45.07" />
                    <SPLIT distance="300" swimtime="00:05:46.99" />
                    <SPLIT distance="350" swimtime="00:06:48.81" />
                    <SPLIT distance="400" swimtime="00:07:50.70" />
                    <SPLIT distance="450" swimtime="00:08:52.25" />
                    <SPLIT distance="500" swimtime="00:09:56.05" />
                    <SPLIT distance="550" swimtime="00:10:57.58" />
                    <SPLIT distance="600" swimtime="00:12:00.52" />
                    <SPLIT distance="650" swimtime="00:13:03.99" />
                    <SPLIT distance="700" swimtime="00:14:06.45" />
                    <SPLIT distance="750" swimtime="00:15:10.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7259" name="MASTERS Zdzieszowice">
          <ATHLETES>
            <ATHLETE firstname="Dorota" lastname="Woźniak" birthdate="1973-09-18" gender="F" nation="POL" swrid="4992846" athleteid="7260">
              <RESULTS>
                <RESULT eventid="1058" points="527" reactiontime="+91" swimtime="00:01:25.45" resultid="7261" heatid="7744" lane="7" entrytime="00:01:25.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="514" reactiontime="+77" swimtime="00:03:03.24" resultid="7262" heatid="7787" lane="6" entrytime="00:03:11.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                    <SPLIT distance="100" swimtime="00:01:29.39" />
                    <SPLIT distance="150" swimtime="00:02:17.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7300" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jarosław" lastname="Tuszyński" birthdate="1975-01-01" gender="M" nation="POL" athleteid="7299">
              <RESULTS>
                <RESULT eventid="1110" points="547" reactiontime="+87" swimtime="00:00:37.03" resultid="7301" heatid="7755" lane="0" entrytime="00:00:36.90" />
                <RESULT eventid="1213" points="312" reactiontime="+93" swimtime="00:00:35.17" resultid="7302" heatid="7770" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1333" points="418" reactiontime="+95" swimtime="00:03:17.39" resultid="7303" heatid="7782" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                    <SPLIT distance="100" swimtime="00:01:35.06" />
                    <SPLIT distance="150" swimtime="00:02:27.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12914" nation="POL" region="14" clubid="7591" name="Water Squad">
          <ATHLETES>
            <ATHLETE firstname="Arkadiusz" lastname="Aptewicz" birthdate="1993-12-20" gender="M" nation="POL" license="112914700053" swrid="4806379" athleteid="7614">
              <RESULTS>
                <RESULT eventid="1110" points="773" reactiontime="+70" swimtime="00:00:30.29" resultid="7615" heatid="7755" lane="6" entrytime="00:00:30.89" entrycourse="SCM" />
                <RESULT eventid="1435" points="856" swimtime="00:08:45.55" resultid="7616" heatid="7792" lane="4" entrytime="00:08:50.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                    <SPLIT distance="100" swimtime="00:01:01.64" />
                    <SPLIT distance="150" swimtime="00:01:34.67" />
                    <SPLIT distance="200" swimtime="00:02:08.11" />
                    <SPLIT distance="250" swimtime="00:02:41.35" />
                    <SPLIT distance="300" swimtime="00:03:14.11" />
                    <SPLIT distance="350" swimtime="00:03:47.24" />
                    <SPLIT distance="400" swimtime="00:04:20.75" />
                    <SPLIT distance="450" swimtime="00:04:54.18" />
                    <SPLIT distance="500" swimtime="00:05:27.84" />
                    <SPLIT distance="550" swimtime="00:06:01.24" />
                    <SPLIT distance="600" swimtime="00:06:34.64" />
                    <SPLIT distance="650" swimtime="00:07:07.92" />
                    <SPLIT distance="700" swimtime="00:07:41.49" />
                    <SPLIT distance="750" swimtime="00:08:14.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Timea" lastname="Balajcza" birthdate="1971-09-22" gender="F" nation="POL" license="512914600062" swrid="5240601" athleteid="7596">
              <RESULTS>
                <RESULT eventid="1058" points="610" reactiontime="+79" swimtime="00:01:21.43" resultid="7597" heatid="7744" lane="3" entrytime="00:01:22.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1093" points="844" reactiontime="+76" swimtime="00:00:37.88" resultid="7598" heatid="7751" lane="3" entrytime="00:00:38.05" entrycourse="SCM" />
                <RESULT eventid="1315" points="722" reactiontime="+81" swimtime="00:03:07.44" resultid="7599" heatid="7779" lane="5" entrytime="00:03:04.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:01:28.44" />
                    <SPLIT distance="150" swimtime="00:02:17.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" license="512914700063" swrid="4655152" athleteid="7603">
              <RESULTS>
                <RESULT eventid="1075" points="198" reactiontime="+80" swimtime="00:01:52.78" resultid="7604" heatid="7746" lane="6" entrytime="00:01:39.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1110" points="369" reactiontime="+83" swimtime="00:00:42.52" resultid="7605" heatid="7754" lane="0" entrytime="00:00:42.48" entrycourse="SCM" />
                <RESULT eventid="1213" points="316" reactiontime="+73" swimtime="00:00:38.19" resultid="7606" heatid="7768" lane="6" entrytime="00:00:37.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Szyszkowska" birthdate="1996-11-05" gender="F" nation="POL" license="512914600054" swrid="4282341" athleteid="7607">
              <RESULTS>
                <RESULT eventid="1093" points="779" swimtime="00:00:34.33" resultid="7608" heatid="7751" lane="4" entrytime="00:00:34.52" entrycourse="SCM" />
                <RESULT eventid="1196" points="766" swimtime="00:00:27.64" resultid="7609" heatid="7766" lane="4" entrytime="00:00:27.66" entrycourse="SCM" />
                <RESULT eventid="1315" points="827" swimtime="00:02:43.71" resultid="7610" heatid="7779" lane="4" entrytime="00:02:40.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                    <SPLIT distance="100" swimtime="00:01:20.38" />
                    <SPLIT distance="150" swimtime="00:02:02.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Kulisz" birthdate="1977-06-16" gender="M" nation="POL" license="512914700002" swrid="5416809" athleteid="7645">
              <RESULTS>
                <RESULT eventid="1145" points="416" reactiontime="+84" swimtime="00:00:34.38" resultid="7646" heatid="7758" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1213" points="508" reactiontime="+90" swimtime="00:00:29.90" resultid="7647" heatid="7771" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1367" reactiontime="+88" status="DNF" swimtime="00:00:00.00" resultid="7648" heatid="7785" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:01:30.90" />
                    <SPLIT distance="150" swimtime="00:02:29.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Kaczmarek" birthdate="1985-05-07" gender="F" nation="POL" license="512914600004" swrid="5240932" athleteid="7592">
              <RESULTS>
                <RESULT eventid="1058" points="797" swimtime="00:01:11.37" resultid="7593" heatid="7744" lane="4" entrytime="00:01:12.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" status="DNS" swimtime="00:00:00.00" resultid="7594" heatid="7762" lane="4" entrytime="00:00:32.42" entrycourse="SCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski w danej kat. wiekowej" eventid="1384" points="812" reactiontime="+78" swimtime="00:02:33.05" resultid="7595" heatid="7787" lane="4" entrytime="00:02:34.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:15.92" />
                    <SPLIT distance="150" swimtime="00:01:55.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Korpetta" birthdate="1959-12-27" gender="M" nation="POL" license="112914700013" swrid="4754654" athleteid="7638">
              <RESULTS>
                <RESULT eventid="1075" points="383" reactiontime="+106" swimtime="00:01:34.01" resultid="7639" heatid="7746" lane="5" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="523" reactiontime="+74" swimtime="00:03:14.90" resultid="7640" heatid="7789" lane="7" entrytime="00:03:15.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                    <SPLIT distance="100" swimtime="00:01:35.45" />
                    <SPLIT distance="150" swimtime="00:02:26.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Dąbrowska" birthdate="1987-05-20" gender="F" nation="POL" license="512914600064" swrid="4655165" athleteid="7621">
              <RESULTS>
                <RESULT eventid="1128" points="213" swimtime="00:00:47.55" resultid="7622" heatid="7757" lane="8" entrytime="00:00:47.35" entrycourse="SCM" />
                <RESULT eventid="1162" points="210" reactiontime="+105" swimtime="00:00:51.96" resultid="7623" heatid="7762" lane="1" entrytime="00:00:52.01" entrycourse="SCM" />
                <RESULT eventid="1196" points="277" swimtime="00:00:40.13" resultid="7624" heatid="7766" lane="9" entrytime="00:00:38.61" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aneta" lastname="Dolińska" birthdate="1990-07-06" gender="F" nation="POL" license="512914600056" swrid="4251116" athleteid="7641">
              <RESULTS>
                <RESULT eventid="1058" points="436" reactiontime="+79" swimtime="00:01:25.49" resultid="7642" heatid="7744" lane="1" entrytime="00:01:26.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="524" swimtime="00:00:32.11" resultid="7643" heatid="7766" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1384" points="371" reactiontime="+84" swimtime="00:03:17.02" resultid="7644" heatid="7787" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                    <SPLIT distance="100" swimtime="00:01:36.79" />
                    <SPLIT distance="150" swimtime="00:02:27.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bożena" lastname="Ayomo" birthdate="1966-02-08" gender="F" nation="POL" license="512914600061" swrid="5582447" athleteid="7600">
              <RESULTS>
                <RESULT eventid="1058" points="389" reactiontime="+90" swimtime="00:01:39.90" resultid="7601" heatid="7743" lane="5" entrytime="00:01:40.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="417" reactiontime="+82" swimtime="00:00:45.28" resultid="7602" heatid="7762" lane="3" entrytime="00:00:44.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Bukowska" birthdate="1985-09-30" gender="F" nation="POL" athleteid="7652">
              <RESULTS>
                <RESULT eventid="1058" points="604" swimtime="00:01:18.29" resultid="7653" heatid="7744" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1093" points="572" reactiontime="+81" swimtime="00:00:38.13" resultid="7654" heatid="7751" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Matyszewski" birthdate="1971-10-11" gender="M" nation="POL" license="512914700065" swrid="5582459" athleteid="7617">
              <RESULTS>
                <RESULT eventid="1110" points="487" reactiontime="+72" swimtime="00:00:39.09" resultid="7618" heatid="7754" lane="5" entrytime="00:00:38.92" entrycourse="SCM" />
                <RESULT eventid="1213" points="373" swimtime="00:00:34.02" resultid="7619" heatid="7769" lane="2" entrytime="00:00:33.83" entrycourse="SCM" />
                <RESULT eventid="1333" points="455" reactiontime="+88" swimtime="00:03:21.16" resultid="7620" heatid="7782" lane="8" entrytime="00:03:21.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                    <SPLIT distance="100" swimtime="00:01:33.73" />
                    <SPLIT distance="150" swimtime="00:02:27.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Markowski" birthdate="1976-01-04" gender="M" nation="POL" license="512914700011" swrid="5471789" athleteid="7627">
              <RESULTS>
                <RESULT eventid="1075" points="560" swimtime="00:01:12.73" resultid="7628" heatid="7748" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="608" reactiontime="+80" swimtime="00:00:30.31" resultid="7629" heatid="7759" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1367" points="525" reactiontime="+85" swimtime="00:02:43.11" resultid="7630" heatid="7785" lane="3" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:01.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Piaściński" birthdate="1976-09-19" gender="M" nation="POL" license="512914700066" athleteid="7631">
              <RESULTS>
                <RESULT eventid="1075" points="590" swimtime="00:01:11.49" resultid="7632" heatid="7747" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="673" reactiontime="+77" swimtime="00:00:31.80" resultid="7633" heatid="7764" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1401" points="565" reactiontime="+81" swimtime="00:02:39.14" resultid="7634" heatid="7789" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:57.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Romuald" lastname="Kozłowski" birthdate="1966-08-13" gender="M" nation="POL" license="512914700012" swrid="5425564" athleteid="7611">
              <RESULTS>
                <RESULT eventid="1110" points="728" reactiontime="+76" swimtime="00:00:33.90" resultid="7612" heatid="7755" lane="1" entrytime="00:00:33.31" entrycourse="SCM" />
                <RESULT eventid="1213" points="803" reactiontime="+81" swimtime="00:00:28.00" resultid="7613" heatid="7771" lane="5" entrytime="00:00:27.94" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Kośmider" birthdate="1966-03-01" gender="M" nation="POL" license="512914700009" swrid="4992964" athleteid="7649">
              <RESULTS>
                <RESULT eventid="1333" points="701" reactiontime="+78" swimtime="00:03:02.36" resultid="7650" heatid="7782" lane="6" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                    <SPLIT distance="100" swimtime="00:01:28.27" />
                    <SPLIT distance="150" swimtime="00:02:15.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="601" swimtime="00:11:01.23" resultid="7651" heatid="7792" lane="9" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:18.81" />
                    <SPLIT distance="150" swimtime="00:02:00.39" />
                    <SPLIT distance="200" swimtime="00:02:42.40" />
                    <SPLIT distance="250" swimtime="00:03:24.94" />
                    <SPLIT distance="300" swimtime="00:04:07.23" />
                    <SPLIT distance="350" swimtime="00:04:49.55" />
                    <SPLIT distance="400" swimtime="00:05:31.77" />
                    <SPLIT distance="450" swimtime="00:06:13.10" />
                    <SPLIT distance="500" swimtime="00:06:54.49" />
                    <SPLIT distance="550" swimtime="00:07:36.21" />
                    <SPLIT distance="600" swimtime="00:08:17.89" />
                    <SPLIT distance="650" swimtime="00:08:59.31" />
                    <SPLIT distance="700" swimtime="00:09:40.30" />
                    <SPLIT distance="750" swimtime="00:10:21.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kaczmarek" birthdate="1977-06-25" gender="M" nation="POL" license="512914700003" swrid="4043251" athleteid="7635">
              <RESULTS>
                <RESULT eventid="1145" points="1029" reactiontime="+72" swimtime="00:00:25.43" resultid="7636" heatid="7760" lane="5" entrytime="00:00:25.15" />
                <RESULT comment="Czas lepszy od Rekordu Polski w danej kat. wiekowej" eventid="1401" points="1002" reactiontime="+72" swimtime="00:02:11.47" resultid="7637" heatid="7789" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:05.11" />
                    <SPLIT distance="150" swimtime="00:01:39.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1247" reactiontime="+79" swimtime="00:05:26.31" resultid="7625" heatid="7774" lane="4" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:10.89" />
                    <SPLIT distance="150" swimtime="00:01:48.49" />
                    <SPLIT distance="200" swimtime="00:02:31.06" />
                    <SPLIT distance="250" swimtime="00:03:07.13" />
                    <SPLIT distance="300" swimtime="00:03:51.17" />
                    <SPLIT distance="350" swimtime="00:04:35.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7631" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="7611" number="2" />
                    <RELAYPOSITION athleteid="7645" number="3" />
                    <RELAYPOSITION athleteid="7603" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski w danej kat. wiekowej" eventid="7052" reactiontime="+67" swimtime="00:05:05.13" resultid="7626" heatid="7775" lane="4" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                    <SPLIT distance="100" swimtime="00:01:30.12" />
                    <SPLIT distance="150" swimtime="00:02:10.90" />
                    <SPLIT distance="200" swimtime="00:02:55.83" />
                    <SPLIT distance="250" swimtime="00:03:22.94" />
                    <SPLIT distance="300" swimtime="00:03:53.55" />
                    <SPLIT distance="350" swimtime="00:04:27.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7638" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="7652" number="2" />
                    <RELAYPOSITION athleteid="7614" number="3" />
                    <RELAYPOSITION athleteid="7641" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7255" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Szymański" birthdate="1978-01-01" gender="M" nation="POL" athleteid="7254">
              <RESULTS>
                <RESULT eventid="1213" points="571" reactiontime="+79" swimtime="00:00:28.76" resultid="7258" heatid="7771" lane="0" entrytime="00:00:29.23" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02805" nation="POL" region="05" clubid="7450" name="MUKS Zgierz">
          <ATHLETES>
            <ATHLETE firstname="Jarosław" lastname="Woźniak" birthdate="1980-09-30" gender="M" nation="POL" license="502805700158" swrid="5506643" athleteid="7498">
              <RESULTS>
                <RESULT eventid="1110" points="364" swimtime="00:00:40.71" resultid="7499" heatid="7754" lane="8" entrytime="00:00:42.18" entrycourse="SCM" />
                <RESULT eventid="1213" points="353" reactiontime="+91" swimtime="00:00:32.82" resultid="7500" heatid="7769" lane="6" entrytime="00:00:33.72" entrycourse="SCM" />
                <RESULT eventid="1333" points="279" reactiontime="+94" swimtime="00:03:38.53" resultid="7501" heatid="7780" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.99" />
                    <SPLIT distance="100" swimtime="00:01:40.22" />
                    <SPLIT distance="150" swimtime="00:02:38.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Matczak" birthdate="1989-08-12" gender="M" nation="POL" license="102805700157" swrid="4071609" athleteid="7492">
              <RESULTS>
                <RESULT eventid="1110" points="802" reactiontime="+69" swimtime="00:00:29.93" resultid="7493" heatid="7755" lane="5" entrytime="00:00:29.77" entrycourse="SCM" />
                <RESULT eventid="1333" points="889" swimtime="00:02:26.13" resultid="7494" heatid="7782" lane="4" entrytime="00:02:21.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:10.17" />
                    <SPLIT distance="150" swimtime="00:01:48.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Ścibiorek" birthdate="1971-09-12" gender="F" nation="POL" license="502805600026" swrid="4992745" athleteid="7470">
              <RESULTS>
                <RESULT eventid="1093" points="810" swimtime="00:00:38.41" resultid="7471" heatid="7751" lane="2" entrytime="00:00:38.92" entrycourse="SCM" />
                <RESULT eventid="1128" points="862" swimtime="00:00:32.72" resultid="7472" heatid="7757" lane="4" entrytime="00:00:32.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Sypniewski" birthdate="1957-02-01" gender="M" nation="POL" license="102805700035" swrid="5373999" athleteid="7451">
              <RESULTS>
                <RESULT eventid="1075" points="587" reactiontime="+76" swimtime="00:01:24.47" resultid="7452" heatid="7747" lane="1" entrytime="00:01:27.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="599" reactiontime="+73" swimtime="00:00:39.52" resultid="7453" heatid="7764" lane="2" entrytime="00:00:40.07" entrycourse="SCM" />
                <RESULT eventid="1333" points="564" reactiontime="+73" swimtime="00:03:39.89" resultid="7454" heatid="7782" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.15" />
                    <SPLIT distance="100" swimtime="00:01:41.36" />
                    <SPLIT distance="150" swimtime="00:02:39.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Rudziński" birthdate="1966-05-10" gender="M" nation="POL" license="502805700162" swrid="4934041" athleteid="7489">
              <RESULTS>
                <RESULT eventid="1110" points="353" reactiontime="+90" swimtime="00:00:43.12" resultid="7490" heatid="7753" lane="5" entrytime="00:00:43.67" entrycourse="SCM" />
                <RESULT eventid="1367" points="224" swimtime="00:03:48.70" resultid="7491" heatid="7784" lane="4" entrytime="00:03:49.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.16" />
                    <SPLIT distance="100" swimtime="00:01:48.05" />
                    <SPLIT distance="150" swimtime="00:02:48.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisław" lastname="Jasiński" birthdate="1960-07-23" gender="M" nation="POL" license="502805700027" swrid="5374015" athleteid="7485">
              <RESULTS>
                <RESULT eventid="1110" points="393" swimtime="00:00:44.68" resultid="7486" heatid="7753" lane="2" entrytime="00:00:44.40" entrycourse="SCM" />
                <RESULT eventid="1213" points="484" reactiontime="+76" swimtime="00:00:34.17" resultid="7487" heatid="7769" lane="7" entrytime="00:00:33.95" entrycourse="SCM" />
                <RESULT eventid="1333" points="397" reactiontime="+98" swimtime="00:03:45.66" resultid="7488" heatid="7781" lane="6" entrytime="00:03:43.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.57" />
                    <SPLIT distance="100" swimtime="00:01:46.81" />
                    <SPLIT distance="150" swimtime="00:02:47.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Klusek" birthdate="1975-01-12" gender="F" nation="POL" license="502805600030" swrid="5464092" athleteid="7473">
              <RESULTS>
                <RESULT eventid="1093" points="561" reactiontime="+88" swimtime="00:00:42.15" resultid="7474" heatid="7749" lane="3" />
                <RESULT eventid="1128" points="526" reactiontime="+93" swimtime="00:00:37.17" resultid="7475" heatid="7756" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Wiśniewska" birthdate="1981-02-26" gender="F" nation="POL" license="502805600123" swrid="5464096" athleteid="7466">
              <RESULTS>
                <RESULT eventid="1093" points="214" reactiontime="+101" swimtime="00:00:57.37" resultid="7467" heatid="7750" lane="6" entrytime="00:00:58.74" entrycourse="SCM" />
                <RESULT eventid="1128" points="120" reactiontime="+112" swimtime="00:00:59.29" resultid="7468" heatid="7757" lane="7" entrytime="00:00:46.20" />
                <RESULT eventid="1196" points="173" reactiontime="+87" swimtime="00:00:47.09" resultid="7469" heatid="7765" lane="5" entrytime="00:00:46.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Pietruszewski - Gil" birthdate="1986-12-17" gender="M" nation="POL" license="502805700163" athleteid="7459">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="7460" heatid="7746" lane="9" />
                <RESULT eventid="1213" points="342" swimtime="00:00:31.50" resultid="7461" heatid="7767" lane="2" />
                <RESULT eventid="1435" status="OTL" swimtime="00:12:07.05" resultid="7793" heatid="7791" lane="9" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="250" swimtime="00:03:32.31" />
                    <SPLIT distance="350" swimtime="00:05:08.73" />
                    <SPLIT distance="400" swimtime="00:09:55.40" />
                    <SPLIT distance="750" swimtime="00:11:27.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Chwiałkowski" birthdate="1985-11-09" gender="M" nation="POL" license="502805700033" swrid="5464089" athleteid="7514">
              <RESULTS>
                <RESULT eventid="1213" points="332" reactiontime="+96" swimtime="00:00:31.81" resultid="7515" heatid="7770" lane="7" entrytime="00:00:31.15" entrycourse="SCM" />
                <RESULT eventid="1435" status="OTL" swimtime="00:12:23.03" resultid="7516" heatid="7791" lane="4" entrytime="00:11:34.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:21.13" />
                    <SPLIT distance="150" swimtime="00:02:05.92" />
                    <SPLIT distance="200" swimtime="00:02:52.16" />
                    <SPLIT distance="250" swimtime="00:03:38.49" />
                    <SPLIT distance="300" swimtime="00:04:25.58" />
                    <SPLIT distance="350" swimtime="00:05:12.52" />
                    <SPLIT distance="400" swimtime="00:06:00.03" />
                    <SPLIT distance="450" swimtime="00:06:48.72" />
                    <SPLIT distance="500" swimtime="00:07:36.28" />
                    <SPLIT distance="550" swimtime="00:08:25.54" />
                    <SPLIT distance="600" swimtime="00:09:14.69" />
                    <SPLIT distance="650" swimtime="00:10:01.85" />
                    <SPLIT distance="700" swimtime="00:10:49.69" />
                    <SPLIT distance="750" swimtime="00:11:37.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Rembowska-Świeboda" birthdate="1968-06-27" gender="F" nation="POL" license="102805600031" swrid="5439505" athleteid="7511">
              <RESULTS>
                <RESULT eventid="1162" points="707" reactiontime="+68" swimtime="00:00:37.98" resultid="7512" heatid="7761" lane="3" />
                <RESULT eventid="1196" points="606" reactiontime="+81" swimtime="00:00:33.94" resultid="7513" heatid="7766" lane="7" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Kajdos" birthdate="1976-06-25" gender="F" nation="POL" license="502805600148" swrid="5558379" athleteid="7508">
              <RESULTS>
                <RESULT eventid="1162" points="249" reactiontime="+110" swimtime="00:00:48.44" resultid="7509" heatid="7762" lane="7" entrytime="00:00:49.96" entrycourse="SCM" />
                <RESULT eventid="1384" points="243" swimtime="00:04:06.39" resultid="7510" heatid="7786" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.24" />
                    <SPLIT distance="100" swimtime="00:03:02.44" />
                    <SPLIT distance="150" swimtime="00:04:06.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Mróz" birthdate="1962-03-03" gender="F" nation="POL" license="502805600024" swrid="4754660" athleteid="7502">
              <RESULTS>
                <RESULT eventid="1128" points="797" reactiontime="+87" swimtime="00:00:36.05" resultid="7503" heatid="7757" lane="3" entrytime="00:00:35.50" entrycourse="SCM" />
                <RESULT eventid="1196" points="735" swimtime="00:00:34.35" resultid="7504" heatid="7766" lane="2" entrytime="00:00:33.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Sikorski" birthdate="1951-05-03" gender="M" nation="POL" license="502805700036" swrid="5582462" athleteid="7495">
              <RESULTS>
                <RESULT eventid="1110" points="278" swimtime="00:00:54.41" resultid="7496" heatid="7753" lane="9" entrytime="00:00:53.03" entrycourse="SCM" />
                <RESULT eventid="1333" points="278" reactiontime="+120" swimtime="00:04:43.60" resultid="7497" heatid="7780" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.61" />
                    <SPLIT distance="100" swimtime="00:02:16.15" />
                    <SPLIT distance="150" swimtime="00:03:32.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tadeusz" lastname="Obiedziński" birthdate="1959-05-12" gender="M" nation="POL" license="502805700040" swrid="4992722" athleteid="7482">
              <RESULTS>
                <RESULT eventid="1110" points="440" swimtime="00:00:43.04" resultid="7483" heatid="7753" lane="4" entrytime="00:00:43.34" entrycourse="SCM" />
                <RESULT eventid="1333" points="310" reactiontime="+96" swimtime="00:04:05.13" resultid="7484" heatid="7781" lane="1" entrytime="00:03:59.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.60" />
                    <SPLIT distance="100" swimtime="00:01:58.22" />
                    <SPLIT distance="150" swimtime="00:03:04.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Morozowski" birthdate="1973-05-09" gender="M" nation="POL" license="102805700051" swrid="5416829" athleteid="7479">
              <RESULTS>
                <RESULT eventid="1110" points="508" reactiontime="+93" swimtime="00:00:38.55" resultid="7480" heatid="7754" lane="6" entrytime="00:00:39.30" entrycourse="SCM" />
                <RESULT eventid="1435" points="344" reactiontime="+112" swimtime="00:12:46.76" resultid="7481" heatid="7791" lane="3" entrytime="00:12:37.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                    <SPLIT distance="100" swimtime="00:01:23.03" />
                    <SPLIT distance="150" swimtime="00:02:08.46" />
                    <SPLIT distance="200" swimtime="00:02:56.29" />
                    <SPLIT distance="250" swimtime="00:03:44.83" />
                    <SPLIT distance="300" swimtime="00:04:34.00" />
                    <SPLIT distance="350" swimtime="00:05:23.52" />
                    <SPLIT distance="400" swimtime="00:06:13.06" />
                    <SPLIT distance="450" swimtime="00:07:04.40" />
                    <SPLIT distance="500" swimtime="00:07:54.54" />
                    <SPLIT distance="550" swimtime="00:08:44.46" />
                    <SPLIT distance="600" swimtime="00:09:34.71" />
                    <SPLIT distance="650" swimtime="00:10:24.50" />
                    <SPLIT distance="700" swimtime="00:11:14.33" />
                    <SPLIT distance="750" swimtime="00:12:02.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="502805600152" swrid="5464091" athleteid="7517">
              <RESULTS>
                <RESULT eventid="1315" points="391" reactiontime="+97" swimtime="00:03:51.47" resultid="7518" heatid="7779" lane="1" entrytime="00:03:50.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.06" />
                    <SPLIT distance="100" swimtime="00:01:50.37" />
                    <SPLIT distance="150" swimtime="00:02:51.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="241" reactiontime="+112" swimtime="00:03:55.10" resultid="7519" heatid="7783" lane="3" entrytime="00:03:53.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.50" />
                    <SPLIT distance="100" swimtime="00:01:52.14" />
                    <SPLIT distance="150" swimtime="00:02:54.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="307" reactiontime="+99" swimtime="00:14:13.12" resultid="7520" heatid="7790" lane="7" entrytime="00:14:05.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.42" />
                    <SPLIT distance="100" swimtime="00:01:40.12" />
                    <SPLIT distance="150" swimtime="00:02:33.95" />
                    <SPLIT distance="200" swimtime="00:03:26.72" />
                    <SPLIT distance="250" swimtime="00:04:19.32" />
                    <SPLIT distance="300" swimtime="00:05:12.62" />
                    <SPLIT distance="350" swimtime="00:06:06.24" />
                    <SPLIT distance="400" swimtime="00:07:00.03" />
                    <SPLIT distance="450" swimtime="00:07:54.26" />
                    <SPLIT distance="500" swimtime="00:08:49.78" />
                    <SPLIT distance="550" swimtime="00:09:44.38" />
                    <SPLIT distance="600" swimtime="00:10:39.54" />
                    <SPLIT distance="650" swimtime="00:11:32.56" />
                    <SPLIT distance="700" swimtime="00:12:27.29" />
                    <SPLIT distance="750" swimtime="00:13:21.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1977-01-05" gender="F" nation="POL" license="502805600055" swrid="4655158" athleteid="7462">
              <RESULTS>
                <RESULT eventid="1093" points="446" reactiontime="+76" swimtime="00:00:45.48" resultid="7463" heatid="7751" lane="1" entrytime="00:00:45.35" entrycourse="SCM" />
                <RESULT eventid="1162" points="275" reactiontime="+86" swimtime="00:00:46.87" resultid="7464" heatid="7762" lane="6" entrytime="00:00:44.40" />
                <RESULT eventid="1315" points="471" swimtime="00:03:37.42" resultid="7465" heatid="7779" lane="6" entrytime="00:03:36.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.15" />
                    <SPLIT distance="100" swimtime="00:01:45.63" />
                    <SPLIT distance="150" swimtime="00:02:42.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Dziedziczak" birthdate="1977-02-04" gender="M" nation="POL" license="502805700153" swrid="5558378" athleteid="7455">
              <RESULTS>
                <RESULT eventid="1075" points="385" swimtime="00:01:22.40" resultid="7456" heatid="7747" lane="2" entrytime="00:01:22.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="385" swimtime="00:00:35.27" resultid="7457" heatid="7758" lane="2" entrytime="00:00:34.46" entrycourse="SCM" />
                <RESULT eventid="1213" points="442" swimtime="00:00:31.32" resultid="7458" heatid="7770" lane="2" entrytime="00:00:31.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Wiczel" birthdate="1948-01-22" gender="M" nation="POL" license="502805700021" swrid="4876444" athleteid="7476">
              <RESULTS>
                <RESULT eventid="1110" points="757" reactiontime="+96" swimtime="00:00:43.00" resultid="7477" heatid="7753" lane="3" entrytime="00:00:44.02" entrycourse="SCM" />
                <RESULT eventid="1333" points="747" reactiontime="+104" swimtime="00:03:35.46" resultid="7478" heatid="7781" lane="3" entrytime="00:03:37.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.22" />
                    <SPLIT distance="100" swimtime="00:01:46.53" />
                    <SPLIT distance="150" swimtime="00:02:42.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dagmara" lastname="Luzniakowska" birthdate="1980-04-29" gender="F" nation="POL" license="102805600154" swrid="5582458" athleteid="7505">
              <RESULTS>
                <RESULT eventid="1128" points="313" swimtime="00:00:43.14" resultid="7506" heatid="7757" lane="2" entrytime="00:00:43.42" entrycourse="SCM" />
                <RESULT eventid="1196" points="372" swimtime="00:00:36.52" resultid="7507" heatid="7765" lane="4" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1247" reactiontime="+80" swimtime="00:05:18.78" resultid="7522" heatid="7774" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                    <SPLIT distance="100" swimtime="00:01:31.54" />
                    <SPLIT distance="150" swimtime="00:02:02.60" />
                    <SPLIT distance="200" swimtime="00:02:37.74" />
                    <SPLIT distance="250" swimtime="00:03:20.36" />
                    <SPLIT distance="300" swimtime="00:04:07.60" />
                    <SPLIT distance="350" swimtime="00:04:40.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7451" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="7492" number="2" />
                    <RELAYPOSITION athleteid="7459" number="3" />
                    <RELAYPOSITION athleteid="7514" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1247" reactiontime="+78" swimtime="00:06:27.67" resultid="7523" heatid="7774" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.92" />
                    <SPLIT distance="100" swimtime="00:01:48.43" />
                    <SPLIT distance="150" swimtime="00:02:37.45" />
                    <SPLIT distance="200" swimtime="00:03:34.67" />
                    <SPLIT distance="250" swimtime="00:04:19.07" />
                    <SPLIT distance="300" swimtime="00:05:14.76" />
                    <SPLIT distance="350" swimtime="00:05:49.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7498" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="7482" number="2" reactiontime="+110" />
                    <RELAYPOSITION athleteid="7489" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="7455" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="7044" reactiontime="+74" swimtime="00:05:35.67" resultid="7521" heatid="7773" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:01:22.99" />
                    <SPLIT distance="150" swimtime="00:02:04.08" />
                    <SPLIT distance="200" swimtime="00:02:50.18" />
                    <SPLIT distance="250" swimtime="00:03:28.78" />
                    <SPLIT distance="300" swimtime="00:04:16.22" />
                    <SPLIT distance="350" swimtime="00:04:54.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7511" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="7470" number="2" />
                    <RELAYPOSITION athleteid="7473" number="3" />
                    <RELAYPOSITION athleteid="7502" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="7052" reactiontime="+100" swimtime="00:06:28.96" resultid="7524" heatid="7775" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.13" />
                    <SPLIT distance="100" swimtime="00:01:50.80" />
                    <SPLIT distance="150" swimtime="00:02:37.96" />
                    <SPLIT distance="200" swimtime="00:03:32.96" />
                    <SPLIT distance="250" swimtime="00:04:13.43" />
                    <SPLIT distance="300" swimtime="00:05:08.41" />
                    <SPLIT distance="350" swimtime="00:05:46.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7508" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="7479" number="2" />
                    <RELAYPOSITION athleteid="7505" number="3" />
                    <RELAYPOSITION athleteid="7485" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7330" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Izabela" lastname="Wypych-Staszewska" birthdate="1970-01-01" gender="F" nation="POL" athleteid="7329">
              <RESULTS>
                <RESULT eventid="1350" points="345" reactiontime="+83" swimtime="00:03:34.17" resultid="7331" heatid="7783" lane="5" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.40" />
                    <SPLIT distance="100" swimtime="00:01:45.79" />
                    <SPLIT distance="150" swimtime="00:02:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="303" reactiontime="+82" swimtime="00:03:38.45" resultid="7332" heatid="7787" lane="8" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.49" />
                    <SPLIT distance="100" swimtime="00:01:46.41" />
                    <SPLIT distance="150" swimtime="00:02:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="358" swimtime="00:13:43.98" resultid="7333" heatid="7790" lane="2" entrytime="00:13:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                    <SPLIT distance="100" swimtime="00:01:33.65" />
                    <SPLIT distance="150" swimtime="00:02:24.98" />
                    <SPLIT distance="200" swimtime="00:03:16.13" />
                    <SPLIT distance="250" swimtime="00:04:07.77" />
                    <SPLIT distance="300" swimtime="00:04:59.96" />
                    <SPLIT distance="350" swimtime="00:05:51.92" />
                    <SPLIT distance="400" swimtime="00:06:44.39" />
                    <SPLIT distance="450" swimtime="00:07:38.06" />
                    <SPLIT distance="500" swimtime="00:08:30.72" />
                    <SPLIT distance="550" swimtime="00:09:23.74" />
                    <SPLIT distance="600" swimtime="00:10:16.83" />
                    <SPLIT distance="650" swimtime="00:11:09.52" />
                    <SPLIT distance="700" swimtime="00:12:02.92" />
                    <SPLIT distance="750" swimtime="00:12:55.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7225" name="Gdynia Masters">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Skwarło" birthdate="1939-01-01" gender="M" nation="POL" swrid="4302086" athleteid="7226">
              <RESULTS>
                <RESULT eventid="1110" points="378" reactiontime="+149" swimtime="00:00:59.45" resultid="7227" heatid="7752" lane="5" entrytime="00:00:57.50" />
                <RESULT eventid="1213" points="170" swimtime="00:00:57.89" resultid="7228" heatid="7767" lane="4" entrytime="00:00:54.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Gorbaczow" birthdate="1987-01-01" gender="M" nation="POL" athleteid="7233">
              <RESULTS>
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /G8" eventid="1075" status="DSQ" swimtime="00:00:00.00" resultid="7234" heatid="7746" lane="4" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="374" reactiontime="+86" swimtime="00:00:30.55" resultid="7235" heatid="7770" lane="8" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Gorbaczow" birthdate="1958-01-01" gender="M" nation="POL" swrid="4191113" athleteid="7229">
              <RESULTS>
                <RESULT eventid="1145" points="870" reactiontime="+79" swimtime="00:00:32.01" resultid="7230" heatid="7758" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1213" points="764" swimtime="00:00:30.16" resultid="7231" heatid="7770" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1401" points="652" reactiontime="+91" swimtime="00:03:01.76" resultid="7232" heatid="7789" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                    <SPLIT distance="100" swimtime="00:01:27.22" />
                    <SPLIT distance="150" swimtime="00:02:15.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7208" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Wiśniewski" birthdate="1973-01-01" gender="M" nation="POL" athleteid="7207">
              <RESULTS>
                <RESULT eventid="1110" points="385" reactiontime="+74" swimtime="00:00:42.25" resultid="7209" heatid="7753" lane="0" entrytime="00:00:51.23" />
                <RESULT eventid="1213" points="391" reactiontime="+70" swimtime="00:00:33.47" resultid="7210" heatid="7769" lane="1" entrytime="00:00:34.27" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7264" name="Weteran Zabrze">
          <ATHLETES>
            <ATHLETE firstname="Krystyna" lastname="Fecica" birthdate="1943-01-01" gender="F" nation="POL" swrid="4102524" athleteid="7263">
              <RESULTS>
                <RESULT eventid="1093" points="676" swimtime="00:00:56.11" resultid="7265" heatid="7750" lane="3" entrytime="00:00:56.00" />
                <RESULT eventid="1128" points="740" swimtime="00:00:53.91" resultid="7266" heatid="7756" lane="4" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7673" name="Swim Club Masters Ślęza">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Chudoba" birthdate="1981-03-04" gender="M" nation="POL" athleteid="7674">
              <RESULTS>
                <RESULT eventid="1075" points="624" reactiontime="+80" swimtime="00:01:10.00" resultid="7675" heatid="7748" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="671" swimtime="00:00:28.70" resultid="7676" heatid="7760" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1367" status="DNS" swimtime="00:00:00.00" resultid="7677" heatid="7785" lane="2" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Sikorski" birthdate="1973-01-18" gender="M" nation="POL" athleteid="7682">
              <RESULTS>
                <RESULT eventid="1110" points="453" swimtime="00:00:40.03" resultid="7683" heatid="7754" lane="2" entrytime="00:00:40.25" />
                <RESULT eventid="1145" points="292" reactiontime="+80" swimtime="00:00:40.39" resultid="7684" heatid="7758" lane="7" entrytime="00:00:39.02" />
                <RESULT eventid="1298" points="365" swimtime="00:00:34.26" resultid="7685" heatid="7777" lane="4" entrytime="00:00:33.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Dusza" birthdate="1983-10-11" gender="F" nation="POL" athleteid="7678">
              <RESULTS>
                <RESULT eventid="1058" points="380" reactiontime="+86" swimtime="00:01:34.06" resultid="7679" heatid="7744" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="355" swimtime="00:00:37.11" resultid="7680" heatid="7766" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1418" points="387" swimtime="00:13:08.68" resultid="7681" heatid="7790" lane="6" entrytime="00:13:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:01:28.76" />
                    <SPLIT distance="150" swimtime="00:02:17.81" />
                    <SPLIT distance="200" swimtime="00:03:07.75" />
                    <SPLIT distance="250" swimtime="00:03:57.57" />
                    <SPLIT distance="300" swimtime="00:04:47.53" />
                    <SPLIT distance="350" swimtime="00:05:37.83" />
                    <SPLIT distance="400" swimtime="00:06:28.43" />
                    <SPLIT distance="450" swimtime="00:07:19.14" />
                    <SPLIT distance="500" swimtime="00:08:09.02" />
                    <SPLIT distance="550" swimtime="00:09:00.17" />
                    <SPLIT distance="600" swimtime="00:09:50.45" />
                    <SPLIT distance="650" swimtime="00:10:40.67" />
                    <SPLIT distance="700" swimtime="00:11:31.53" />
                    <SPLIT distance="750" swimtime="00:12:21.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7221" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Bołtuć" birthdate="1983-01-01" gender="F" nation="POL" athleteid="7220">
              <RESULTS>
                <RESULT eventid="1058" points="395" swimtime="00:01:32.81" resultid="7222" heatid="7743" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="401" reactiontime="+126" swimtime="00:03:22.59" resultid="7223" heatid="7787" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.60" />
                    <SPLIT distance="100" swimtime="00:01:41.23" />
                    <SPLIT distance="150" swimtime="00:02:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="509" reactiontime="+102" swimtime="00:11:59.91" resultid="7224" heatid="7790" lane="5" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:24.11" />
                    <SPLIT distance="150" swimtime="00:02:09.03" />
                    <SPLIT distance="200" swimtime="00:02:54.55" />
                    <SPLIT distance="250" swimtime="00:03:40.28" />
                    <SPLIT distance="300" swimtime="00:04:25.46" />
                    <SPLIT distance="350" swimtime="00:05:11.03" />
                    <SPLIT distance="400" swimtime="00:05:57.05" />
                    <SPLIT distance="450" swimtime="00:06:43.03" />
                    <SPLIT distance="500" swimtime="00:07:28.51" />
                    <SPLIT distance="550" swimtime="00:08:14.12" />
                    <SPLIT distance="600" swimtime="00:08:59.80" />
                    <SPLIT distance="650" swimtime="00:09:45.35" />
                    <SPLIT distance="700" swimtime="00:10:30.38" />
                    <SPLIT distance="750" swimtime="00:11:16.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TMBAR" nation="POL" clubid="7124" name="Tm Barracuda">
          <ATHLETES>
            <ATHLETE firstname="Karolina" lastname="Stasiak" birthdate="1984-05-06" gender="F" nation="POL" license="505815600033" athleteid="7129">
              <RESULTS>
                <RESULT eventid="1093" points="266" reactiontime="+96" swimtime="00:00:49.20" resultid="7130" heatid="7751" lane="0" entrytime="00:00:49.61" />
                <RESULT eventid="1128" points="206" reactiontime="+91" swimtime="00:00:48.13" resultid="7131" heatid="7757" lane="0" entrytime="00:00:48.34" />
                <RESULT eventid="1315" points="337" swimtime="00:03:42.83" resultid="7132" heatid="7779" lane="2" entrytime="00:03:43.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.35" />
                    <SPLIT distance="100" swimtime="00:01:47.04" />
                    <SPLIT distance="150" swimtime="00:02:44.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Radomska" birthdate="1982-04-12" gender="F" nation="POL" license="505815600016" athleteid="7125">
              <RESULTS>
                <RESULT eventid="1058" points="361" swimtime="00:01:35.66" resultid="7126" heatid="7744" lane="9" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="436" reactiontime="+82" swimtime="00:00:34.65" resultid="7127" heatid="7766" lane="1" entrytime="00:00:34.72" />
                <RESULT eventid="1418" points="390" reactiontime="+94" swimtime="00:13:06.57" resultid="7128" heatid="7790" lane="3" entrytime="00:13:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                    <SPLIT distance="100" swimtime="00:01:26.34" />
                    <SPLIT distance="150" swimtime="00:02:13.91" />
                    <SPLIT distance="200" swimtime="00:03:02.49" />
                    <SPLIT distance="250" swimtime="00:03:53.16" />
                    <SPLIT distance="300" swimtime="00:04:42.31" />
                    <SPLIT distance="350" swimtime="00:05:33.89" />
                    <SPLIT distance="400" swimtime="00:06:23.90" />
                    <SPLIT distance="450" swimtime="00:07:14.81" />
                    <SPLIT distance="500" swimtime="00:08:05.27" />
                    <SPLIT distance="550" swimtime="00:08:56.56" />
                    <SPLIT distance="600" swimtime="00:09:46.91" />
                    <SPLIT distance="650" swimtime="00:10:37.44" />
                    <SPLIT distance="700" swimtime="00:11:27.98" />
                    <SPLIT distance="750" swimtime="00:12:18.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="GBR" clubid="7077" name="Cardiff">
          <ATHLETES>
            <ATHLETE firstname="Marco" lastname="Menegazzi" birthdate="1980-01-01" gender="M" nation="GBR" athleteid="7076">
              <RESULTS>
                <RESULT eventid="1145" points="566" swimtime="00:00:30.38" resultid="7078" heatid="7759" lane="2" entrytime="00:00:30.29" />
                <RESULT eventid="1213" points="527" reactiontime="+83" swimtime="00:00:28.73" resultid="7079" heatid="7771" lane="1" entrytime="00:00:28.52" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="7106" name="Ukraine Swim Team">
          <ATHLETES>
            <ATHLETE firstname="Natalia" lastname="Boryshkevych" birthdate="1976-04-15" gender="F" nation="UKR" swrid="5241793" athleteid="7105">
              <RESULTS>
                <RESULT eventid="1058" points="642" reactiontime="+65" swimtime="00:01:20.10" resultid="7107" heatid="7744" lane="6" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="628" swimtime="00:11:12.28" resultid="7108" heatid="7790" lane="4" entrytime="00:11:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                    <SPLIT distance="150" swimtime="00:02:00.53" />
                    <SPLIT distance="200" swimtime="00:02:43.07" />
                    <SPLIT distance="250" swimtime="00:03:25.71" />
                    <SPLIT distance="300" swimtime="00:04:08.50" />
                    <SPLIT distance="350" swimtime="00:04:51.47" />
                    <SPLIT distance="400" swimtime="00:05:34.66" />
                    <SPLIT distance="450" swimtime="00:06:18.09" />
                    <SPLIT distance="500" swimtime="00:07:01.53" />
                    <SPLIT distance="550" swimtime="00:07:44.60" />
                    <SPLIT distance="600" swimtime="00:08:27.67" />
                    <SPLIT distance="650" swimtime="00:09:09.82" />
                    <SPLIT distance="700" swimtime="00:09:51.85" />
                    <SPLIT distance="750" swimtime="00:10:33.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02016" nation="POL" region="16" clubid="7370" name="Koszalińskie TKKF">
          <ATHLETES>
            <ATHLETE firstname="Grzegorz" lastname="Ćwikła" birthdate="1974-08-22" gender="M" nation="POL" license="102016700002" swrid="5506628" athleteid="7377">
              <RESULTS>
                <RESULT eventid="1179" points="573" reactiontime="+75" swimtime="00:00:33.54" resultid="7378" heatid="7764" lane="6" entrytime="00:00:33.36" entrycourse="SCM" />
                <RESULT eventid="1401" points="515" swimtime="00:02:44.10" resultid="7379" heatid="7789" lane="5" entrytime="00:02:44.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="150" swimtime="00:02:01.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="436" reactiontime="+89" swimtime="00:11:25.19" resultid="7380" heatid="7792" lane="8" entrytime="00:10:52.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                    <SPLIT distance="100" swimtime="00:01:17.55" />
                    <SPLIT distance="150" swimtime="00:01:59.82" />
                    <SPLIT distance="200" swimtime="00:02:42.60" />
                    <SPLIT distance="250" swimtime="00:03:25.49" />
                    <SPLIT distance="300" swimtime="00:04:08.96" />
                    <SPLIT distance="350" swimtime="00:04:52.36" />
                    <SPLIT distance="400" swimtime="00:05:35.84" />
                    <SPLIT distance="450" swimtime="00:06:19.71" />
                    <SPLIT distance="500" swimtime="00:07:03.92" />
                    <SPLIT distance="550" swimtime="00:07:48.02" />
                    <SPLIT distance="600" swimtime="00:08:32.48" />
                    <SPLIT distance="650" swimtime="00:09:16.36" />
                    <SPLIT distance="700" swimtime="00:10:00.36" />
                    <SPLIT distance="750" swimtime="00:10:43.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Rutkowski" birthdate="1951-10-06" gender="M" nation="POL" license="102016700022" swrid="5506639" athleteid="7371">
              <RESULTS>
                <RESULT eventid="1075" points="265" swimtime="00:02:00.75" resultid="7372" heatid="7746" lane="2" entrytime="00:01:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="283" swimtime="00:00:43.24" resultid="7373" heatid="7768" lane="8" entrytime="00:00:43.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Rutkowski" birthdate="1974-02-20" gender="M" nation="POL" license="102016700018" swrid="4992794" athleteid="7374">
              <RESULTS>
                <RESULT eventid="1145" points="550" reactiontime="+77" swimtime="00:00:31.33" resultid="7375" heatid="7759" lane="1" entrytime="00:00:31.80" />
                <RESULT eventid="1367" points="413" reactiontime="+84" swimtime="00:02:56.68" resultid="7376" heatid="7785" lane="7" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:21.30" />
                    <SPLIT distance="150" swimtime="00:02:08.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="7560" name="Warsaw Masters Team">
          <ATHLETES>
            <ATHLETE firstname="Dymitr" lastname="Bielski" birthdate="1977-08-13" gender="M" nation="POL" license="104214700039" swrid="5552366" athleteid="7564">
              <RESULTS>
                <RESULT eventid="1075" points="471" reactiontime="+94" swimtime="00:01:17.05" resultid="7565" heatid="7747" lane="6" entrytime="00:01:17.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="459" reactiontime="+81" swimtime="00:00:30.94" resultid="7566" heatid="7770" lane="5" entrytime="00:00:30.80" entrycourse="SCM" />
                <RESULT eventid="1435" points="438" reactiontime="+92" swimtime="00:11:24.28" resultid="7567" heatid="7792" lane="0" entrytime="00:11:18.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:16.96" />
                    <SPLIT distance="150" swimtime="00:01:58.16" />
                    <SPLIT distance="200" swimtime="00:02:40.08" />
                    <SPLIT distance="250" swimtime="00:03:23.41" />
                    <SPLIT distance="350" swimtime="00:05:34.87" />
                    <SPLIT distance="500" swimtime="00:07:01.27" />
                    <SPLIT distance="550" swimtime="00:07:44.90" />
                    <SPLIT distance="600" swimtime="00:08:29.87" />
                    <SPLIT distance="650" swimtime="00:09:13.55" />
                    <SPLIT distance="700" swimtime="00:09:58.13" />
                    <SPLIT distance="750" swimtime="00:10:41.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Szemberg" birthdate="1949-07-26" gender="F" nation="POL" license="504214600017" swrid="4302692" athleteid="7561">
              <RESULTS>
                <RESULT eventid="1058" points="159" swimtime="00:02:33.86" resultid="7562" heatid="7743" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="397" swimtime="00:17:45.62" resultid="7563" heatid="7790" lane="8" entrytime="00:18:08.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.89" />
                    <SPLIT distance="100" swimtime="00:02:06.84" />
                    <SPLIT distance="150" swimtime="00:03:15.49" />
                    <SPLIT distance="200" swimtime="00:04:22.45" />
                    <SPLIT distance="250" swimtime="00:05:29.83" />
                    <SPLIT distance="300" swimtime="00:06:37.15" />
                    <SPLIT distance="350" swimtime="00:07:43.74" />
                    <SPLIT distance="400" swimtime="00:08:49.74" />
                    <SPLIT distance="450" swimtime="00:09:57.71" />
                    <SPLIT distance="500" swimtime="00:11:04.83" />
                    <SPLIT distance="550" swimtime="00:12:12.13" />
                    <SPLIT distance="600" swimtime="00:13:18.83" />
                    <SPLIT distance="650" swimtime="00:14:24.89" />
                    <SPLIT distance="700" swimtime="00:15:32.09" />
                    <SPLIT distance="750" swimtime="00:16:38.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Warchoł" birthdate="1953-08-30" gender="M" nation="POL" license="504214700035" swrid="4222718" athleteid="7584">
              <RESULTS>
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /G8" eventid="1075" status="DSQ" swimtime="00:00:00.00" resultid="7585" heatid="7745" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="1197" reactiontime="+107" swimtime="00:02:51.35" resultid="7586" heatid="7788" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:22.52" />
                    <SPLIT distance="150" swimtime="00:02:08.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Skośkiewicz" birthdate="1966-05-05" gender="M" nation="POL" license="504214700002" swrid="4183802" athleteid="7572">
              <RESULTS>
                <RESULT eventid="1075" points="910" reactiontime="+77" swimtime="00:01:07.82" resultid="7573" heatid="7748" lane="6" entrytime="00:01:10.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="780" swimtime="00:00:30.46" resultid="7574" heatid="7759" lane="4" entrytime="00:00:29.92" entrycourse="SCM" />
                <RESULT eventid="1401" points="811" reactiontime="+71" swimtime="00:02:33.55" resultid="7575" heatid="7788" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:55.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leszek" lastname="Madej" birthdate="1960-06-17" gender="M" nation="POL" license="504214700005" swrid="4183799" athleteid="7568">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="7569" heatid="7748" lane="8" entrytime="00:01:11.11" entrycourse="SCM" />
                <RESULT eventid="1145" status="DNS" swimtime="00:00:00.00" resultid="7570" heatid="7759" lane="9" entrytime="00:00:32.17" entrycourse="SCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="7571" heatid="7771" lane="4" entrytime="00:00:27.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Rogosz" birthdate="1976-04-28" gender="M" nation="POL" license="504214700003" swrid="4270348" athleteid="7576">
              <RESULTS>
                <RESULT eventid="1075" points="579" reactiontime="+86" swimtime="00:01:11.94" resultid="7577" heatid="7745" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="556" reactiontime="+87" swimtime="00:00:29.02" resultid="7578" heatid="7767" lane="3" />
                <RESULT eventid="1435" points="567" reactiontime="+102" swimtime="00:10:27.97" resultid="7579" heatid="7792" lane="7" entrytime="00:10:44.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:01:13.67" />
                    <SPLIT distance="150" swimtime="00:01:53.45" />
                    <SPLIT distance="200" swimtime="00:02:33.72" />
                    <SPLIT distance="250" swimtime="00:03:13.79" />
                    <SPLIT distance="300" swimtime="00:03:53.84" />
                    <SPLIT distance="350" swimtime="00:04:33.61" />
                    <SPLIT distance="400" swimtime="00:05:13.25" />
                    <SPLIT distance="450" swimtime="00:05:52.83" />
                    <SPLIT distance="500" swimtime="00:06:32.32" />
                    <SPLIT distance="550" swimtime="00:07:12.51" />
                    <SPLIT distance="600" swimtime="00:07:52.36" />
                    <SPLIT distance="650" swimtime="00:08:32.15" />
                    <SPLIT distance="700" swimtime="00:09:12.18" />
                    <SPLIT distance="750" swimtime="00:09:51.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Paluszak" birthdate="1967-02-17" gender="M" nation="POL" license="504214700102" swrid="5471792" athleteid="7580">
              <RESULTS>
                <RESULT eventid="1075" points="305" swimtime="00:01:37.64" resultid="7581" heatid="7746" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="283" swimtime="00:00:42.70" resultid="7582" heatid="7758" lane="9" />
                <RESULT eventid="1213" points="274" swimtime="00:00:40.04" resultid="7583" heatid="7767" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ostrowski" birthdate="1977-05-14" gender="M" nation="POL" license="504214700091" swrid="5506635" athleteid="7587">
              <RESULTS>
                <RESULT eventid="1110" points="913" swimtime="00:00:31.22" resultid="7588" heatid="7755" lane="2" entrytime="00:00:31.89" entrycourse="SCM" />
                <RESULT eventid="1333" points="692" reactiontime="+76" swimtime="00:02:46.92" resultid="7589" heatid="7782" lane="3" entrytime="00:02:48.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:16.57" />
                    <SPLIT distance="150" swimtime="00:02:02.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="529" reactiontime="+78" swimtime="00:10:42.72" resultid="7590" heatid="7792" lane="1" entrytime="00:10:45.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:13.86" />
                    <SPLIT distance="150" swimtime="00:01:53.69" />
                    <SPLIT distance="200" swimtime="00:02:34.36" />
                    <SPLIT distance="250" swimtime="00:03:14.82" />
                    <SPLIT distance="300" swimtime="00:03:55.41" />
                    <SPLIT distance="350" swimtime="00:04:36.09" />
                    <SPLIT distance="400" swimtime="00:05:17.01" />
                    <SPLIT distance="450" swimtime="00:05:58.53" />
                    <SPLIT distance="500" swimtime="00:06:40.08" />
                    <SPLIT distance="550" swimtime="00:07:20.95" />
                    <SPLIT distance="600" swimtime="00:08:01.98" />
                    <SPLIT distance="650" swimtime="00:08:42.79" />
                    <SPLIT distance="700" swimtime="00:09:23.95" />
                    <SPLIT distance="750" swimtime="00:10:04.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" nation="POL" clubid="7133" name="KS Masters Polkowice">
          <ATHLETES>
            <ATHLETE firstname="Emilia" lastname="Kawula" birthdate="1941-10-02" gender="F" nation="POL" athleteid="7158">
              <RESULTS>
                <RESULT eventid="1093" points="40" swimtime="00:02:23.48" resultid="7159" heatid="7749" lane="4" entrytime="00:02:17.00" entrycourse="SCM" />
                <RESULT eventid="1196" points="110" swimtime="00:01:27.81" resultid="7160" heatid="7765" lane="7" entrytime="00:01:33.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogdan" lastname="Jawor" birthdate="1947-04-23" gender="M" nation="POL" swrid="4754745" athleteid="7134">
              <RESULTS>
                <RESULT eventid="1075" points="289" reactiontime="+90" swimtime="00:02:06.34" resultid="7135" heatid="7746" lane="7" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="205" reactiontime="+98" swimtime="00:01:01.71" resultid="7136" heatid="7763" lane="6" entrytime="00:01:01.00" entrycourse="SCM" />
                <RESULT eventid="1401" points="232" reactiontime="+135" swimtime="00:04:52.85" resultid="7137" heatid="7788" lane="6" entrytime="00:04:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.33" />
                    <SPLIT distance="100" swimtime="00:02:21.34" />
                    <SPLIT distance="150" swimtime="00:03:38.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kazimierz" lastname="Rosik" birthdate="1955-11-11" gender="M" nation="POL" athleteid="7146">
              <RESULTS>
                <RESULT eventid="1110" points="301" swimtime="00:00:50.40" resultid="7147" heatid="7752" lane="4" entrytime="00:00:54.00" entrycourse="SCM" />
                <RESULT eventid="1213" points="265" reactiontime="+106" swimtime="00:00:42.91" resultid="7148" heatid="7768" lane="0" entrytime="00:00:44.00" entrycourse="SCM" />
                <RESULT eventid="1333" points="388" reactiontime="+120" swimtime="00:04:08.99" resultid="7149" heatid="7781" lane="8" entrytime="00:04:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.37" />
                    <SPLIT distance="100" swimtime="00:01:58.73" />
                    <SPLIT distance="150" swimtime="00:03:03.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Świder" birthdate="1943-11-28" gender="F" nation="POL" athleteid="7161">
              <RESULTS>
                <RESULT eventid="1093" points="81" swimtime="00:01:53.48" resultid="7162" heatid="7750" lane="1" entrytime="00:01:38.00" entrycourse="SCM" />
                <RESULT eventid="1196" points="109" swimtime="00:01:28.03" resultid="7163" heatid="7765" lane="1" entrytime="00:01:39.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiesław" lastname="Zając" birthdate="1946-01-02" gender="M" nation="POL" athleteid="7142">
              <RESULTS>
                <RESULT eventid="1110" points="165" reactiontime="+106" swimtime="00:01:11.47" resultid="7143" heatid="7752" lane="3" entrytime="00:01:13.00" entrycourse="SCM" />
                <RESULT eventid="1179" points="95" reactiontime="+97" swimtime="00:01:19.54" resultid="7144" heatid="7763" lane="2" entrytime="00:01:14.00" entrycourse="SCM" />
                <RESULT eventid="1333" points="196" reactiontime="+106" swimtime="00:05:36.31" resultid="7145" heatid="7781" lane="0" entrytime="00:05:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.94" />
                    <SPLIT distance="100" swimtime="00:02:43.01" />
                    <SPLIT distance="150" swimtime="00:04:15.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisława" lastname="Pachom" birthdate="1945-10-10" gender="F" nation="POL" athleteid="7154">
              <RESULTS>
                <RESULT eventid="1093" points="59" swimtime="00:02:00.87" resultid="7155" heatid="7750" lane="8" entrytime="00:01:50.00" entrycourse="SCM" />
                <RESULT eventid="1162" points="64" swimtime="00:01:48.90" resultid="7156" heatid="7761" lane="5" entrytime="00:01:50.00" entrycourse="SCM" />
                <RESULT eventid="1196" points="59" swimtime="00:01:28.37" resultid="7157" heatid="7765" lane="2" entrytime="00:01:33.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gizela" lastname="Wójcik" birthdate="1949-11-16" gender="F" nation="POL" athleteid="7175">
              <RESULTS>
                <RESULT eventid="1093" points="215" swimtime="00:01:12.00" resultid="7176" heatid="7750" lane="7" entrytime="00:01:15.00" entrycourse="SCM" />
                <RESULT eventid="1162" points="227" reactiontime="+162" swimtime="00:01:08.49" resultid="7177" heatid="7762" lane="8" entrytime="00:01:10.00" entrycourse="SCM" />
                <RESULT eventid="1315" points="272" swimtime="00:05:29.07" resultid="7178" heatid="7778" lane="6" entrytime="00:05:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.11" />
                    <SPLIT distance="100" swimtime="00:02:38.47" />
                    <SPLIT distance="150" swimtime="00:04:03.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Regina" lastname="Mładszew" birthdate="1952-07-15" gender="F" nation="POL" athleteid="7150">
              <RESULTS>
                <RESULT eventid="1058" points="101" reactiontime="+123" swimtime="00:02:58.57" resultid="7151" heatid="7743" lane="7" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="147" reactiontime="+187" swimtime="00:01:19.19" resultid="7152" heatid="7761" lane="4" entrytime="00:01:29.00" entrycourse="SCM" />
                <RESULT eventid="1384" points="163" reactiontime="+143" swimtime="00:06:01.60" resultid="7153" heatid="7787" lane="0" entrytime="00:05:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.19" />
                    <SPLIT distance="100" swimtime="00:03:01.30" />
                    <SPLIT distance="150" swimtime="00:04:33.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Ołpiński" birthdate="1991-04-26" gender="M" nation="POL" swrid="4217107" athleteid="7164">
              <RESULTS>
                <RESULT eventid="1145" points="483" reactiontime="+77" swimtime="00:00:29.13" resultid="7165" heatid="7760" lane="0" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1213" points="504" swimtime="00:00:27.80" resultid="7166" heatid="7772" lane="9" entrytime="00:00:27.25" entrycourse="SCM" />
                <RESULT eventid="1333" points="351" swimtime="00:03:19.17" resultid="7167" heatid="7782" lane="2" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                    <SPLIT distance="100" swimtime="00:01:32.81" />
                    <SPLIT distance="150" swimtime="00:02:26.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Leśniak" birthdate="1957-03-27" gender="F" nation="POL" athleteid="7168">
              <RESULTS>
                <RESULT eventid="1196" points="50" swimtime="00:01:27.12" resultid="7169" heatid="7765" lane="6" entrytime="00:01:30.00" entrycourse="SCM" />
                <RESULT eventid="1384" points="88" swimtime="00:07:03.44" resultid="7170" heatid="7786" lane="4" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.78" />
                    <SPLIT distance="100" swimtime="00:03:33.63" />
                    <SPLIT distance="150" swimtime="00:05:18.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janina" lastname="Zając" birthdate="1946-08-16" gender="F" nation="POL" athleteid="7138">
              <RESULTS>
                <RESULT eventid="1093" points="138" swimtime="00:01:31.08" resultid="7139" heatid="7750" lane="0" entrytime="00:01:53.80" entrycourse="SCM" />
                <RESULT eventid="1196" points="116" swimtime="00:01:10.77" resultid="7140" heatid="7765" lane="3" entrytime="00:01:11.00" entrycourse="SCM" />
                <RESULT eventid="1384" points="163" reactiontime="+56" swimtime="00:06:10.39" resultid="7141" heatid="7786" lane="5" entrytime="00:06:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.33" />
                    <SPLIT distance="100" swimtime="00:03:01.25" />
                    <SPLIT distance="150" swimtime="00:04:37.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zygmunt" lastname="Pawlaczek" birthdate="1949-05-26" gender="M" nation="POL" athleteid="7171">
              <RESULTS>
                <RESULT eventid="1110" points="379" reactiontime="+101" swimtime="00:00:49.08" resultid="7172" heatid="7753" lane="1" entrytime="00:00:48.60" entrycourse="SCM" />
                <RESULT eventid="1213" points="391" swimtime="00:00:38.83" resultid="7173" heatid="7768" lane="2" entrytime="00:00:38.80" entrycourse="SCM" />
                <RESULT eventid="1435" points="337" reactiontime="+153" swimtime="00:16:27.73" resultid="7174" heatid="7791" lane="8" entrytime="00:16:21.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.39" />
                    <SPLIT distance="100" swimtime="00:01:48.94" />
                    <SPLIT distance="150" swimtime="00:02:46.57" />
                    <SPLIT distance="200" swimtime="00:03:48.42" />
                    <SPLIT distance="250" swimtime="00:04:52.11" />
                    <SPLIT distance="300" swimtime="00:05:56.06" />
                    <SPLIT distance="350" swimtime="00:06:59.19" />
                    <SPLIT distance="400" swimtime="00:08:02.18" />
                    <SPLIT distance="450" swimtime="00:09:06.36" />
                    <SPLIT distance="500" swimtime="00:10:10.47" />
                    <SPLIT distance="550" swimtime="00:11:14.93" />
                    <SPLIT distance="600" swimtime="00:12:20.05" />
                    <SPLIT distance="650" swimtime="00:13:23.73" />
                    <SPLIT distance="700" swimtime="00:14:28.29" />
                    <SPLIT distance="750" swimtime="00:15:30.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORONA 191" nation="POL" clubid="7184" name="Korona1919 Kraków">
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Leńczowska" birthdate="1982-01-15" gender="F" nation="POL" swrid="4992907" athleteid="7192">
              <RESULTS>
                <RESULT eventid="1128" points="602" reactiontime="+80" swimtime="00:00:34.70" resultid="7193" heatid="7757" lane="5" entrytime="00:00:33.70" />
                <RESULT eventid="1162" points="535" reactiontime="+72" swimtime="00:00:37.61" resultid="7194" heatid="7762" lane="5" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Macierzewska" birthdate="1960-04-20" gender="F" nation="POL" swrid="4992827" athleteid="7189">
              <RESULTS>
                <RESULT eventid="1058" points="643" swimtime="00:01:31.63" resultid="7190" heatid="7744" lane="8" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="946" swimtime="00:03:27.01" resultid="7191" heatid="7783" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                    <SPLIT distance="100" swimtime="00:01:36.63" />
                    <SPLIT distance="150" swimtime="00:02:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="603" reactiontime="+89" swimtime="00:00:42.97" resultid="7687" heatid="7762" lane="2" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariola" lastname="Kuliś" birthdate="1966-07-27" gender="F" nation="POL" swrid="4992797" athleteid="7185">
              <RESULTS>
                <RESULT eventid="1093" points="998" reactiontime="+71" swimtime="00:00:37.58" resultid="7186" heatid="7751" lane="6" entrytime="00:00:38.25" />
                <RESULT eventid="1196" points="837" reactiontime="+74" swimtime="00:00:30.48" resultid="7187" heatid="7766" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1384" points="687" reactiontime="+66" swimtime="00:02:57.93" resultid="7188" heatid="7787" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                    <SPLIT distance="100" swimtime="00:01:25.27" />
                    <SPLIT distance="150" swimtime="00:02:11.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Janeczko" birthdate="1972-12-23" gender="F" nation="POL" swrid="4218717" athleteid="7195">
              <RESULTS>
                <RESULT eventid="1058" points="410" reactiontime="+92" swimtime="00:01:32.93" resultid="7196" heatid="7743" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="619" swimtime="00:00:36.54" resultid="7197" heatid="7757" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1384" points="343" reactiontime="+96" swimtime="00:03:29.70" resultid="7198" heatid="7787" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.24" />
                    <SPLIT distance="100" swimtime="00:01:43.61" />
                    <SPLIT distance="150" swimtime="00:02:38.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7211" name="Motyl Mosir Stalowa Wola">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Petecka" birthdate="1967-04-17" gender="F" nation="POL" license="100908600388" swrid="4992840" athleteid="7212">
              <RESULTS>
                <RESULT eventid="1093" points="497" swimtime="00:00:47.40" resultid="7213" heatid="7751" lane="8" entrytime="00:00:49.00" />
                <RESULT eventid="1196" points="475" reactiontime="+85" swimtime="00:00:36.82" resultid="7214" heatid="7766" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1315" points="587" reactiontime="+88" swimtime="00:03:41.24" resultid="7215" heatid="7779" lane="7" entrytime="00:03:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.79" />
                    <SPLIT distance="100" swimtime="00:01:46.05" />
                    <SPLIT distance="150" swimtime="00:02:43.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7343" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Dominik" lastname="Rudzki" birthdate="1992-01-01" gender="M" nation="POL" swrid="4250678" athleteid="7342">
              <RESULTS>
                <RESULT eventid="1075" points="633" swimtime="00:01:04.04" resultid="7344" heatid="7748" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="575" reactiontime="+60" swimtime="00:00:27.49" resultid="7345" heatid="7760" lane="6" entrytime="00:00:27.29" />
                <RESULT eventid="1213" points="633" reactiontime="+60" swimtime="00:00:25.77" resultid="7346" heatid="7772" lane="3" entrytime="00:00:25.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7119" name="MKS Juvenia Białystok">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Żmiejko" birthdate="1963-01-16" gender="M" nation="POL" license="500309700377" swrid="4186249" athleteid="7120">
              <RESULTS>
                <RESULT eventid="1075" points="866" reactiontime="+74" swimtime="00:01:11.62" resultid="7121" heatid="7746" lane="1" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" status="DNS" swimtime="00:00:00.00" resultid="7122" heatid="7759" lane="7" entrytime="00:00:30.67" entrycourse="SCM" />
                <RESULT eventid="1213" points="837" swimtime="00:00:28.48" resultid="7123" heatid="7771" lane="2" entrytime="00:00:28.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00612" nation="POL" region="12" clubid="7385" name="KS KSZO Ostrowiec Św.">
          <ATHLETES>
            <ATHLETE firstname="Stanisław" lastname="Sejmicki" birthdate="1961-05-04" gender="M" nation="POL" license="500612700426" swrid="5558380" athleteid="7386">
              <RESULTS>
                <RESULT eventid="1110" points="480" reactiontime="+96" swimtime="00:00:41.79" resultid="7387" heatid="7753" lane="6" entrytime="00:00:44.35" entrycourse="SCM" />
                <RESULT eventid="1213" points="411" reactiontime="+106" swimtime="00:00:36.08" resultid="7388" heatid="7768" lane="5" entrytime="00:00:36.38" entrycourse="SCM" />
                <RESULT eventid="1333" points="436" swimtime="00:03:38.68" resultid="7389" heatid="7781" lane="2" entrytime="00:03:44.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                    <SPLIT distance="100" swimtime="00:01:43.38" />
                    <SPLIT distance="150" swimtime="00:02:41.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7666" name="Niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Roman" lastname="Domagała" birthdate="2003-01-01" gender="M" nation="POL" swrid="4840761" athleteid="7669">
              <RESULTS>
                <RESULT eventid="1110" points="802" swimtime="00:00:30.41" resultid="7670" heatid="7755" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1213" points="809" swimtime="00:00:24.61" resultid="7671" heatid="7772" lane="4" entrytime="00:00:24.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KTP" nation="POL" clubid="7267" name="Kościańskie Towarzystwo Pływackie">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Pelec" birthdate="1987-01-29" gender="M" nation="POL" athleteid="7278">
              <RESULTS>
                <RESULT eventid="1110" points="198" swimtime="00:00:49.47" resultid="7279" heatid="7754" lane="9" entrytime="00:00:43.00" entrycourse="SCM" />
                <RESULT eventid="1213" points="257" swimtime="00:00:34.65" resultid="7280" heatid="7769" lane="3" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1333" points="210" swimtime="00:03:56.51" resultid="7281" heatid="7781" lane="7" entrytime="00:03:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.52" />
                    <SPLIT distance="100" swimtime="00:01:53.78" />
                    <SPLIT distance="150" swimtime="00:02:55.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Brygier" birthdate="1979-09-05" gender="F" nation="POL" athleteid="7286">
              <RESULTS>
                <RESULT eventid="1058" points="215" swimtime="00:01:53.63" resultid="7287" heatid="7743" lane="2" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="169" reactiontime="+106" swimtime="00:00:52.99" resultid="7288" heatid="7757" lane="1" entrytime="00:00:47.00" entrycourse="SCM" />
                <RESULT eventid="1315" points="278" reactiontime="+120" swimtime="00:04:14.41" resultid="7289" heatid="7778" lane="5" entrytime="00:04:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.58" />
                    <SPLIT distance="100" swimtime="00:02:05.71" />
                    <SPLIT distance="150" swimtime="00:03:11.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Naglik" birthdate="1968-10-27" gender="M" nation="POL" athleteid="7274">
              <RESULTS>
                <RESULT eventid="1179" points="192" reactiontime="+83" swimtime="00:00:50.81" resultid="7275" heatid="7763" lane="5" entrytime="00:00:50.00" entrycourse="SCM" />
                <RESULT eventid="1367" points="178" reactiontime="+99" swimtime="00:04:06.87" resultid="7276" heatid="7784" lane="5" entrytime="00:03:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.94" />
                    <SPLIT distance="100" swimtime="00:01:55.77" />
                    <SPLIT distance="150" swimtime="00:03:02.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="204" reactiontime="+111" swimtime="00:04:03.32" resultid="7277" heatid="7788" lane="5" entrytime="00:03:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.76" />
                    <SPLIT distance="100" swimtime="00:01:59.31" />
                    <SPLIT distance="150" swimtime="00:03:02.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Rychlik" birthdate="1968-03-17" gender="M" nation="POL" athleteid="7268">
              <RESULTS>
                <RESULT eventid="1298" points="19" swimtime="00:01:36.82" resultid="7269" heatid="7777" lane="6" entrytime="00:01:50.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Morawski" birthdate="1991-02-22" gender="M" nation="POL" athleteid="7282">
              <RESULTS>
                <RESULT eventid="1075" points="254" swimtime="00:01:26.83" resultid="7283" heatid="7747" lane="8" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="324" swimtime="00:00:32.19" resultid="7284" heatid="7770" lane="9" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1333" points="299" swimtime="00:03:30.04" resultid="7285" heatid="7782" lane="9" entrytime="00:03:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.38" />
                    <SPLIT distance="100" swimtime="00:01:41.62" />
                    <SPLIT distance="150" swimtime="00:02:34.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewelina" lastname="Braun" birthdate="1976-11-30" gender="F" nation="POL" athleteid="7290">
              <RESULTS>
                <RESULT eventid="1093" points="270" reactiontime="+87" swimtime="00:00:53.75" resultid="7291" heatid="7750" lane="5" entrytime="00:00:55.00" entrycourse="SCM" />
                <RESULT eventid="1315" points="276" swimtime="00:04:19.88" resultid="7292" heatid="7779" lane="8" entrytime="00:03:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.71" />
                    <SPLIT distance="100" swimtime="00:02:00.40" />
                    <SPLIT distance="150" swimtime="00:03:10.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Skrzypczak" birthdate="1966-09-14" gender="M" nation="POL" swrid="4992721" athleteid="7270">
              <RESULTS>
                <RESULT eventid="1179" points="254" reactiontime="+91" swimtime="00:00:46.31" resultid="7271" heatid="7764" lane="0" entrytime="00:00:47.00" entrycourse="SCM" />
                <RESULT eventid="1367" points="304" reactiontime="+92" swimtime="00:03:26.75" resultid="7272" heatid="7785" lane="8" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                    <SPLIT distance="100" swimtime="00:01:37.79" />
                    <SPLIT distance="150" swimtime="00:02:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="294" reactiontime="+88" swimtime="00:03:35.35" resultid="7273" heatid="7789" lane="0" entrytime="00:03:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                    <SPLIT distance="100" swimtime="00:01:45.69" />
                    <SPLIT distance="150" swimtime="00:02:41.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="7052" reactiontime="+88" swimtime="00:07:03.73" resultid="7293" heatid="7775" lane="6" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                    <SPLIT distance="100" swimtime="00:01:39.82" />
                    <SPLIT distance="150" swimtime="00:02:35.67" />
                    <SPLIT distance="200" swimtime="00:03:37.84" />
                    <SPLIT distance="250" swimtime="00:04:29.31" />
                    <SPLIT distance="300" swimtime="00:05:29.86" />
                    <SPLIT distance="350" swimtime="00:06:14.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7270" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="7290" number="2" reactiontime="+71" />
                    <RELAYPOSITION athleteid="7274" number="3" />
                    <RELAYPOSITION athleteid="7286" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7180" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Kęsik" birthdate="1979-01-01" gender="M" nation="POL" athleteid="7179">
              <RESULTS>
                <RESULT eventid="1075" points="798" reactiontime="+71" swimtime="00:01:04.48" resultid="7181" heatid="7748" lane="5" entrytime="00:01:06.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="735" swimtime="00:00:27.84" resultid="7182" heatid="7760" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1213" points="711" swimtime="00:00:26.00" resultid="7183" heatid="7772" lane="2" entrytime="00:00:26.12" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7335" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Klimkowski" birthdate="1981-01-01" gender="M" nation="POL" swrid="4629756" athleteid="7334">
              <RESULTS>
                <RESULT eventid="1179" points="30" swimtime="00:01:26.47" resultid="7336" heatid="7763" lane="7" entrytime="00:01:34.48" />
                <RESULT eventid="1213" points="13" swimtime="00:01:37.73" resultid="7337" heatid="7767" lane="5" entrytime="00:01:36.22" />
                <RESULT eventid="1298" points="13" swimtime="00:01:36.32" resultid="7338" heatid="7777" lane="3" entrytime="00:01:36.22" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10414" nation="POL" region="14" clubid="7358" name="Klub Sportowy Mako">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Kosiela" birthdate="1985-02-03" gender="M" nation="POL" license="510414700076" athleteid="7363">
              <RESULTS>
                <RESULT eventid="1075" points="233" reactiontime="+89" swimtime="00:01:32.18" resultid="7364" heatid="7745" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="235" reactiontime="+96" swimtime="00:00:35.68" resultid="7365" heatid="7767" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Ostapczuk" birthdate="1970-07-13" gender="M" nation="POL" license="510414700077" athleteid="7359">
              <RESULTS>
                <RESULT eventid="1075" points="272" reactiontime="+100" swimtime="00:01:31.45" resultid="7360" heatid="7745" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1110" points="322" reactiontime="+92" swimtime="00:00:44.86" resultid="7361" heatid="7752" lane="6" />
                <RESULT eventid="1213" points="335" reactiontime="+92" swimtime="00:00:35.25" resultid="7362" heatid="7767" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Piórkowski" birthdate="1965-07-28" gender="M" nation="POL" license="510414700072" swrid="5506637" athleteid="7366">
              <RESULTS>
                <RESULT eventid="1179" points="218" reactiontime="+78" swimtime="00:00:48.72" resultid="7367" heatid="7764" lane="9" entrytime="00:00:47.37" entrycourse="SCM" />
                <RESULT eventid="1213" points="299" reactiontime="+91" swimtime="00:00:38.92" resultid="7368" heatid="7768" lane="7" entrytime="00:00:39.56" entrycourse="SCM" />
                <RESULT eventid="1401" points="223" reactiontime="+97" swimtime="00:03:55.99" resultid="7369" heatid="7789" lane="9" entrytime="00:03:43.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.45" />
                    <SPLIT distance="100" swimtime="00:01:57.03" />
                    <SPLIT distance="150" swimtime="00:02:57.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7313" name="UMKSN Poznań">
          <ATHLETES>
            <ATHLETE firstname="Bohdana" lastname="Davydova" birthdate="2004-01-01" gender="F" nation="POL" athleteid="7317">
              <RESULTS>
                <RESULT eventid="7068" points="347" reactiontime="+93" swimtime="00:00:37.01" resultid="7318" heatid="7776" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gordian" lastname="Wypchał" birthdate="2015-01-01" gender="M" nation="POL" athleteid="7327">
              <RESULTS>
                <RESULT eventid="1298" swimtime="00:01:26.65" resultid="7328" heatid="7777" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Borys" lastname="Rozumek" birthdate="2015-01-01" gender="M" nation="POL" athleteid="7325">
              <RESULTS>
                <RESULT eventid="1298" swimtime="00:01:21.58" resultid="7326" heatid="7777" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kornel" lastname="Jarosz" birthdate="2015-01-01" gender="M" nation="POL" athleteid="7323">
              <RESULTS>
                <RESULT eventid="1298" swimtime="00:01:33.19" resultid="7324" heatid="7777" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Lewandowski" birthdate="2003-01-01" gender="M" nation="POL" athleteid="7321">
              <RESULTS>
                <RESULT eventid="1298" points="68" swimtime="00:00:56.18" resultid="7322" heatid="7777" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sandra" lastname="Michałowska" birthdate="1993-01-01" gender="F" nation="POL" swrid="4660596" athleteid="7312">
              <RESULTS>
                <RESULT eventid="7068" points="504" swimtime="00:00:32.54" resultid="7314" heatid="7776" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Kniaź" birthdate="1996-01-01" gender="F" nation="POL" swrid="4258684" athleteid="7315">
              <RESULTS>
                <RESULT eventid="7068" points="231" reactiontime="+114" swimtime="00:00:41.16" resultid="7316" heatid="7776" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Musiał" birthdate="2010-01-01" gender="F" nation="POL" athleteid="7319">
              <RESULTS>
                <RESULT eventid="7068" reactiontime="+101" swimtime="00:00:59.04" resultid="7320" heatid="7776" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" region="11" clubid="7381" name="KS Górnik Radlin">
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Kubica" birthdate="1972-02-22" gender="M" nation="POL" license="100211700343" swrid="5398297" athleteid="7382">
              <RESULTS>
                <RESULT eventid="1145" points="550" swimtime="00:00:32.72" resultid="7383" heatid="7758" lane="4" entrytime="00:00:32.19" entrycourse="SCM" />
                <RESULT eventid="1401" points="496" reactiontime="+81" swimtime="00:02:55.75" resultid="7384" heatid="7789" lane="6" entrytime="00:02:52.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:01:24.94" />
                    <SPLIT distance="150" swimtime="00:02:10.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7236" name="5 Styl Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Barnasiuk" birthdate="1992-02-04" gender="M" nation="POL" swrid="4273597" athleteid="7241">
              <RESULTS>
                <RESULT eventid="1145" points="535" reactiontime="+62" swimtime="00:00:28.17" resultid="7242" heatid="7760" lane="1" entrytime="00:00:28.70" entrycourse="SCM" />
                <RESULT eventid="1213" points="620" reactiontime="+65" swimtime="00:00:25.95" resultid="7243" heatid="7772" lane="1" entrytime="00:00:27.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Niedzwiadek" birthdate="1993-10-18" gender="M" nation="POL" athleteid="7244">
              <RESULTS>
                <RESULT eventid="1213" points="476" reactiontime="+83" swimtime="00:00:28.33" resultid="7245" heatid="7771" lane="7" entrytime="00:00:28.20" entrycourse="SCM" />
                <RESULT eventid="1435" points="642" reactiontime="+74" swimtime="00:09:38.52" resultid="7246" heatid="7792" lane="5" entrytime="00:09:38.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:43.29" />
                    <SPLIT distance="200" swimtime="00:02:19.91" />
                    <SPLIT distance="250" swimtime="00:02:56.19" />
                    <SPLIT distance="300" swimtime="00:03:33.07" />
                    <SPLIT distance="350" swimtime="00:04:09.76" />
                    <SPLIT distance="400" swimtime="00:04:46.63" />
                    <SPLIT distance="450" swimtime="00:05:23.22" />
                    <SPLIT distance="500" swimtime="00:05:59.71" />
                    <SPLIT distance="550" swimtime="00:06:36.98" />
                    <SPLIT distance="600" swimtime="00:07:13.72" />
                    <SPLIT distance="650" swimtime="00:07:50.22" />
                    <SPLIT distance="700" swimtime="00:08:26.90" />
                    <SPLIT distance="750" swimtime="00:09:04.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Broniszewski" birthdate="1980-09-26" gender="M" nation="POL" athleteid="7237">
              <RESULTS>
                <RESULT eventid="1075" points="325" reactiontime="+80" swimtime="00:01:27.00" resultid="7238" heatid="7747" lane="7" entrytime="00:01:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1110" points="355" reactiontime="+81" swimtime="00:00:41.06" resultid="7239" heatid="7754" lane="3" entrytime="00:00:39.00" entrycourse="SCM" />
                <RESULT eventid="1213" points="336" reactiontime="+80" swimtime="00:00:33.37" resultid="7240" heatid="7769" lane="5" entrytime="00:00:33.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Wziątek" birthdate="1988-01-14" gender="M" nation="POL" athleteid="7247">
              <RESULTS>
                <RESULT eventid="1145" points="340" reactiontime="+78" swimtime="00:00:33.85" resultid="7248" heatid="7759" lane="0" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1435" points="400" reactiontime="+78" swimtime="00:11:36.17" resultid="7249" heatid="7791" lane="5" entrytime="00:12:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                    <SPLIT distance="150" swimtime="00:01:57.58" />
                    <SPLIT distance="200" swimtime="00:02:40.54" />
                    <SPLIT distance="250" swimtime="00:03:24.52" />
                    <SPLIT distance="300" swimtime="00:04:08.41" />
                    <SPLIT distance="350" swimtime="00:04:52.51" />
                    <SPLIT distance="400" swimtime="00:05:37.15" />
                    <SPLIT distance="450" swimtime="00:06:22.65" />
                    <SPLIT distance="500" swimtime="00:07:07.90" />
                    <SPLIT distance="550" swimtime="00:07:53.35" />
                    <SPLIT distance="600" swimtime="00:08:38.85" />
                    <SPLIT distance="650" swimtime="00:09:23.90" />
                    <SPLIT distance="700" swimtime="00:10:09.32" />
                    <SPLIT distance="750" swimtime="00:10:54.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1247" reactiontime="+78" swimtime="00:04:59.49" resultid="7250" heatid="7774" lane="5" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="150" swimtime="00:01:50.23" />
                    <SPLIT distance="200" swimtime="00:02:37.97" />
                    <SPLIT distance="250" swimtime="00:03:12.93" />
                    <SPLIT distance="300" swimtime="00:03:57.19" />
                    <SPLIT distance="350" swimtime="00:04:26.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7241" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="7237" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="7247" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="7244" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02706" nation="POL" region="06" clubid="7534" name="UKS ,,Jasień&apos;&apos; Sucha Beskidzka">
          <ATHLETES>
            <ATHLETE firstname="Sabina" lastname="Sikora" birthdate="1984-10-03" gender="F" nation="POL" license="102706600159" swrid="5468086" athleteid="7535">
              <RESULTS>
                <RESULT eventid="1093" points="677" reactiontime="+73" swimtime="00:00:36.05" resultid="7536" heatid="7751" lane="5" entrytime="00:00:35.13" entrycourse="SCM" />
                <RESULT eventid="1196" points="659" reactiontime="+71" swimtime="00:00:30.07" resultid="7537" heatid="7766" lane="5" entrytime="00:00:29.28" entrycourse="SCM" />
                <RESULT eventid="1315" points="584" reactiontime="+73" swimtime="00:03:05.53" resultid="7538" heatid="7779" lane="3" entrytime="00:03:05.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:01:30.20" />
                    <SPLIT distance="150" swimtime="00:02:18.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7662" name="Niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Sokulski" birthdate="1991-01-01" gender="M" nation="POL" swrid="4062177" athleteid="7661">
              <RESULTS>
                <RESULT eventid="1145" points="725" swimtime="00:00:25.45" resultid="7663" heatid="7760" lane="4" entrytime="00:00:25.00" />
                <RESULT eventid="1213" points="760" reactiontime="+66" swimtime="00:00:24.25" resultid="7664" heatid="7772" lane="5" entrytime="00:00:24.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7309" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Poloch" birthdate="1983-01-01" gender="M" nation="POL" athleteid="7308">
              <RESULTS>
                <RESULT eventid="1110" points="264" reactiontime="+87" swimtime="00:00:45.28" resultid="7310" heatid="7754" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1213" points="366" reactiontime="+88" swimtime="00:00:32.43" resultid="7311" heatid="7769" lane="8" entrytime="00:00:34.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" clubid="7095" name="Ks Extreme Team Oborniki">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Wolniewicz" birthdate="1948-12-22" gender="M" nation="POL" swrid="4754624" athleteid="7096">
              <RESULTS>
                <RESULT eventid="1145" points="232" reactiontime="+104" swimtime="00:00:55.27" resultid="7097" heatid="7758" lane="0" entrytime="00:00:52.00" />
                <RESULT eventid="1213" points="511" reactiontime="+103" swimtime="00:00:39.14" resultid="7098" heatid="7768" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1435" points="330" reactiontime="+113" swimtime="00:17:34.30" resultid="7099" heatid="7791" lane="0" entrytime="00:18:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.30" />
                    <SPLIT distance="100" swimtime="00:01:53.64" />
                    <SPLIT distance="150" swimtime="00:02:57.86" />
                    <SPLIT distance="200" swimtime="00:04:01.92" />
                    <SPLIT distance="250" swimtime="00:05:08.36" />
                    <SPLIT distance="300" swimtime="00:06:15.85" />
                    <SPLIT distance="350" swimtime="00:07:22.83" />
                    <SPLIT distance="400" swimtime="00:08:30.45" />
                    <SPLIT distance="450" swimtime="00:09:38.88" />
                    <SPLIT distance="500" swimtime="00:10:46.70" />
                    <SPLIT distance="550" swimtime="00:11:54.70" />
                    <SPLIT distance="600" swimtime="00:13:03.48" />
                    <SPLIT distance="650" swimtime="00:14:10.87" />
                    <SPLIT distance="700" swimtime="00:15:21.22" />
                    <SPLIT distance="750" swimtime="00:16:29.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01012" nation="POL" region="12" clubid="7445" name="MOSiR Ostrowiec Św.">
          <ATHLETES>
            <ATHLETE firstname="Józef" lastname="Różalski" birthdate="1945-03-28" gender="M" nation="POL" license="501012700001" swrid="4216999" athleteid="7446">
              <RESULTS>
                <RESULT eventid="1110" points="330" reactiontime="+96" swimtime="00:00:56.70" resultid="7447" heatid="7752" lane="7" />
                <RESULT eventid="1213" points="365" swimtime="00:00:43.76" resultid="7448" heatid="7767" lane="6" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="7449" heatid="7780" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7110" name="niezrzeszony Jarocin">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Marszałek" birthdate="1954-10-24" gender="M" nation="POL" athleteid="7109">
              <RESULTS>
                <RESULT eventid="1145" points="179" swimtime="00:00:54.22" resultid="7111" heatid="7758" lane="8" entrytime="00:00:50.40" />
                <RESULT eventid="1213" points="268" reactiontime="+76" swimtime="00:00:42.75" resultid="7112" heatid="7768" lane="1" entrytime="00:00:40.20" />
                <RESULT eventid="1435" points="311" swimtime="00:15:31.47" resultid="7113" heatid="7791" lane="2" entrytime="00:14:44.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.33" />
                    <SPLIT distance="100" swimtime="00:01:51.58" />
                    <SPLIT distance="150" swimtime="00:02:49.94" />
                    <SPLIT distance="200" swimtime="00:03:48.67" />
                    <SPLIT distance="250" swimtime="00:04:47.94" />
                    <SPLIT distance="300" swimtime="00:05:45.99" />
                    <SPLIT distance="350" swimtime="00:06:44.86" />
                    <SPLIT distance="400" swimtime="00:07:43.01" />
                    <SPLIT distance="450" swimtime="00:08:41.97" />
                    <SPLIT distance="500" swimtime="00:09:40.97" />
                    <SPLIT distance="550" swimtime="00:10:39.48" />
                    <SPLIT distance="600" swimtime="00:11:38.12" />
                    <SPLIT distance="650" swimtime="00:12:36.76" />
                    <SPLIT distance="700" swimtime="00:13:35.66" />
                    <SPLIT distance="750" swimtime="00:14:34.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7115" name="niezrzeszony Środa Wlkp.">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Grzelczak" birthdate="1985-10-10" gender="M" nation="POL" athleteid="7114">
              <RESULTS>
                <RESULT eventid="1075" points="200" reactiontime="+100" swimtime="00:01:37.11" resultid="7116" heatid="7746" lane="3" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1110" points="325" reactiontime="+95" swimtime="00:00:41.96" resultid="7117" heatid="7754" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="1333" points="299" swimtime="00:03:30.22" resultid="7118" heatid="7781" lane="4" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.42" />
                    <SPLIT distance="100" swimtime="00:01:38.86" />
                    <SPLIT distance="150" swimtime="00:02:34.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7340" name="niezrzeszony Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Franciszek" lastname="Stasieńko" birthdate="2006-01-01" gender="M" nation="POL" athleteid="7339">
              <RESULTS>
                <RESULT eventid="1298" swimtime="00:00:42.58" resultid="7341" heatid="7777" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03210" nation="POL" region="10" clubid="7435" name="MKP Gdańsk">
          <ATHLETES>
            <ATHLETE firstname="Michalina" lastname="Majewski" birthdate="1984-12-26" gender="F" nation="POL" license="103210600112" athleteid="7436">
              <RESULTS>
                <RESULT eventid="1058" points="691" reactiontime="+79" swimtime="00:01:14.83" resultid="7437" heatid="7743" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1093" points="507" reactiontime="+77" swimtime="00:00:39.69" resultid="7438" heatid="7749" lane="5" />
                <RESULT eventid="1315" points="583" swimtime="00:03:05.68" resultid="7439" heatid="7778" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                    <SPLIT distance="100" swimtime="00:01:30.59" />
                    <SPLIT distance="150" swimtime="00:02:18.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
